VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO an41
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 18.500 BY 30.000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    USE SIGNAL ;
    PORT
      LAYER ML2 ;
        POLYGON 1.000 15.500  1.000 17.500  3.000 17.500  3.000 15.500  1.000 
        15.500  ;
    END
    PORT
      LAYER ML1 ;
        POLYGON 1.000 15.500  1.000 17.500  3.000 17.500  3.000 15.500  1.000 
        15.500  ;
    END
  END A
  PIN B
    USE SIGNAL ;
    PORT
      LAYER ML2 ;
        POLYGON 4.000 12.500  4.000 14.500  6.000 14.500  6.000 12.500  4.000 
        12.500  ;
    END
    PORT
      LAYER ML1 ;
        POLYGON 4.000 12.500  4.000 14.500  6.000 14.500  6.000 12.500  4.000 
        12.500  ;
    END
  END B
  PIN C
    USE SIGNAL ;
    PORT
      LAYER ML2 ;
        POLYGON 7.000 9.700  7.000 11.700  9.000 11.700  9.000 9.700  7.000 
        9.700  ;
    END
    PORT
      LAYER ML1 ;
        POLYGON 7.000 9.700  7.000 11.700  9.000 11.700  9.000 9.700  7.000 
        9.700  ;
    END
  END C
  PIN D
    USE SIGNAL ;
    PORT
      LAYER ML2 ;
        POLYGON 10.000 12.500  10.000 14.500  12.000 14.500  12.000 12.500  
        10.000 12.500  ;
    END
    PORT
      LAYER ML1 ;
        POLYGON 10.000 12.500  10.000 14.500  12.000 14.500  12.000 12.500  
        10.000 12.500  ;
    END
  END D
  PIN VDD
    USE POWER ;
    PORT
      LAYER ML1 ;
        RECT -0.500 28.500  19.000 30.500  ;
    END
  END VDD
  PIN VSS
    USE GROUND ;
    PORT
      LAYER ML1 ;
        RECT -0.500 -0.500  19.000 1.500  ;
    END
  END VSS
  PIN Y
    USE SIGNAL ;
    PORT
      LAYER ML1 ;
        POLYGON 16.000 12.700  16.000 14.700  18.000 14.700  18.000 12.700  
        16.000 12.700  ;
    END
    PORT
      LAYER ML2 ;
        POLYGON 16.000 12.700  16.000 14.700  18.000 14.700  18.000 12.700  
        16.000 12.700  ;
    END
    PORT
      LAYER ML1 ;
        WIDTH 1.000  ;
        PATH 16.800 20.500 16.800 8.000 13.800 8.000 13.800 3.800  ;
    END
  END Y
  OBS
    LAYER ML1 ;
      WIDTH 1.400  ;
      PATH 1.800 21.300 1.800 28.500  ;
      WIDTH 1.000  ;
      PATH 1.800 1.000 1.800 3.800  ;
      WIDTH 1.400  ;
      PATH 4.800 21.300 4.800 24.500  ;
      WIDTH 1.400  ;
      PATH 7.800 21.300 7.800 28.500  ;
      WIDTH 1.000  ;
      PATH 4.800 20.500 4.800 18.000 13.800 18.000 13.800 10.000 10.800 10.000 
      10.800 3.800  ;
      WIDTH 1.000  ;
      PATH 10.800 20.500 10.800 18.000  ;
      WIDTH 1.400  ;
      PATH 10.800 21.300 10.800 24.500  ;
      WIDTH 1.400  ;
      PATH 13.800 21.300 13.800 28.500  ;
      WIDTH 1.400  ;
      PATH 13.800 21.300 13.800 24.500  ;
      WIDTH 1.400  ;
      PATH 16.800 21.300 16.800 24.500  ;
    VIA 1.800 22.500  dcont ;
    VIA 1.800 20.500  dcont ;
    VIA 1.800 3.800  dcont ;
    VIA 1.800 24.500  dcont ;
    VIA 4.800 22.500  dcont ;
    VIA 4.800 20.500  dcont ;
    VIA 4.800 24.500  dcont ;
    VIA 7.800 24.500  dcont ;
    VIA 7.800 22.500  dcont ;
    VIA 7.800 20.500  dcont ;
    VIA 10.800 3.800  dcont ;
    VIA 10.800 20.500  dcont ;
    VIA 10.800 22.500  dcont ;
    VIA 10.800 24.500  dcont ;
    VIA 13.800 24.500  dcont ;
    VIA 13.800 22.500  dcont ;
    VIA 13.800 20.500  dcont ;
    VIA 13.800 3.800  dcont ;
    VIA 16.800 20.500  dcont ;
    VIA 16.800 22.500  dcont ;
    VIA 16.800 24.500  dcont ;
    VIA 14.300 10.500  pcont ;
    VIA 11.000 13.500  pcont ;
    VIA 8.000 10.700  pcont ;
    VIA 5.500 29.500  nsubcont ;
    VIA 5.000 13.500  pcont ;
    VIA 2.000 16.500  pcont ;
    VIA 5.000 0.500  psubcont ;
  END
END an41

MACRO dcont
  CLASS CORE ;
  OBS
    LAYER ML1 ;
      RECT -1.000 -1.000  1.000 1.000  ;
  END
END dcont

MACRO pcont
  CLASS CORE ;
  OBS
    LAYER ML1 ;
      RECT -1.000 -1.000  1.000 1.000  ;
  END
END pcont

MACRO nsubcont
  CLASS CORE ;
  OBS
    LAYER ML1 ;
      RECT -1.000 -1.000  1.000 1.000  ;
  END
END nsubcont

MACRO psubcont
  CLASS CORE ;
  OBS
    LAYER ML1 ;
      RECT -1.000 -1.000  1.000 1.000  ;
  END
END psubcont


END LIBRARY
