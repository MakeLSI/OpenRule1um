VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO or21
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 12.500 BY 30.000 ;
  SYMMETRY X Y ;
  SITE unit ;
 
  PIN A
    USE SIGNAL ;
    PORT
      LAYER ML1 ;
        POLYGON 1.000 8.500  1.000 10.500  3.000 10.500  3.000 8.500  1.000 
        8.500  ;
    END
    PORT
      LAYER ML2 ;
        POLYGON 1.000 8.500  1.000 10.500  3.000 10.500  3.000 8.500  1.000 
        8.500  ;
    END
  END A
  PIN B
    USE SIGNAL ;
    PORT
      LAYER ML1 ;
        POLYGON 4.000 11.500  4.000 13.500  6.000 13.500  6.000 11.500  4.000 
        11.500  ;
    END
    PORT
      LAYER ML2 ;
        POLYGON 4.000 11.500  4.000 13.500  6.000 13.500  6.000 11.500  4.000 
        11.500  ;
    END
  END B
  PIN VDD
    USE POWER ;
    PORT
      LAYER ML1 ;
        RECT -0.500 28.500  13.000 30.500  ;
    END
  END VDD
  PIN VSS
    USE GROUND ;
    PORT
      LAYER ML1 ;
        RECT -0.500 -0.500  13.000 1.500  ;
    END
  END VSS
  PIN Y
    USE SIGNAL ;
    PORT
      LAYER ML1 ;
        WIDTH 1.000  ;
        PATH 10.800 3.800 10.800 18.000 10.300 18.000 10.300 20.500  ;
    END
    PORT
      LAYER ML1 ;
        POLYGON 10.000 8.000  10.000 10.000  12.000 10.000  12.000 8.000  
        10.000 8.000  ;
    END
    PORT
      LAYER ML2 ;
        POLYGON 10.000 8.000  10.000 10.000  12.000 10.000  12.000 8.000  
        10.000 8.000  ;
    END
  END Y
  OBS

    LAYER ML1 ;
      WIDTH 1.000  ;
      PATH 1.800 1.000 1.800 3.800  ;

      WIDTH 1.400  ;
      PATH 2.300 21.300 2.300 24.500  ;

      WIDTH 1.000  ;
      PATH 4.800 3.800 4.800 6.300 7.800 6.300 7.800 16.500 2.300 16.500 2.300 
      20.500  ;

      WIDTH 1.400  ;
      PATH 7.300 21.300 7.300 28.500  ;
      WIDTH 1.000  ;
      PATH 7.800 1.000 7.800 3.800  ;
      WIDTH 1.400  ;
      PATH 10.300 21.300 10.300 24.500  ;
      WIDTH 1.000  ;
      PATH 10.800 3.800 10.800 18.000 10.300 18.000 10.300 20.500  ;

    VIA 1.800 3.800  dcont ;
    VIA 2.300 22.500  dcont ;
    VIA 2.300 20.500  dcont ;
    VIA 2.300 24.500  dcont ;
    VIA 4.800 3.800  dcont ;
    VIA 7.300 20.500  dcont ;
    VIA 7.300 22.500  dcont ;
    VIA 7.300 24.500  dcont ;
    VIA 7.800 3.800  dcont ;
    VIA 10.300 22.500  dcont ;
    VIA 10.300 20.500  dcont ;
    VIA 10.300 24.500  dcont ;
    VIA 10.800 3.800  dcont ;
    VIA 5.500 29.500  nsubcont ;
    VIA 5.000 12.500  pcont ;
    VIA 8.300 12.500  pcont ;
    VIA 2.000 9.500  pcont ;
    VIA 5.000 0.500  psubcont ;
  END
END or21

MACRO dcont
  CLASS CORE ;
  OBS
    LAYER ML1 ;
      RECT -1.000 -1.000  1.000 1.000  ;
  END
END dcont

MACRO nsubcont
  CLASS CORE ;
  OBS
    LAYER ML1 ;
      RECT -1.000 -1.000  1.000 1.000  ;
  END
END nsubcont

MACRO pcont
  CLASS CORE ;
  OBS
    LAYER ML1 ;
      RECT -1.000 -1.000  1.000 1.000  ;
  END
END pcont

MACRO psubcont
  CLASS CORE ;
  OBS
    LAYER ML1 ;
      RECT -1.000 -1.000  1.000 1.000  ;
  END
END psubcont


END LIBRARY
