VERSION 5.3 ;

NAMESCASESENSITIVE ON ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS











MACRO an31
  CLASS BLOCK ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER ML1 ;
        POLYGON 1.000 9.700  1.000 11.700  3.000 11.700  3.000 9.700  1.000 
        9.700  ;
    END
    PORT
      LAYER ML2 ;
        POLYGON 1.000 9.700  1.000 11.700  3.000 11.700  3.000 9.700  1.000 
        9.700  ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER ML1 ;
        POLYGON 4.000 12.500  4.000 14.500  6.000 14.500  6.000 12.500  4.000 
        12.500  ;
    END
    PORT
      LAYER ML2 ;
        POLYGON 4.000 12.500  4.000 14.500  6.000 14.500  6.000 12.500  4.000 
        12.500  ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER ML2 ;
        POLYGON 7.000 9.700  7.000 11.700  9.000 11.700  9.000 9.700  7.000 
        9.700  ;
    END
    PORT
      LAYER ML1 ;
        POLYGON 7.000 9.700  7.000 11.700  9.000 11.700  9.000 9.700  7.000 
        9.700  ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    PORT
      LAYER ML1 ;
        RECT -0.500 28.500  16.000 30.500  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    PORT
      LAYER ML1 ;
        RECT -0.500 -0.500  16.000 1.500  ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    PORT
      LAYER ML2 ;
        POLYGON 13.000 12.700  13.000 14.700  15.000 14.700  15.000 12.700  
        13.000 12.700  ;
    END
    PORT
      LAYER ML1 ;
        POLYGON 13.000 12.700  13.000 14.700  15.000 14.700  15.000 12.700  
        13.000 12.700  ;
    END
    PORT
      LAYER ML1 ;
        WIDTH 1.000  ;
        PATH 13.800 20.500 13.800 3.800 11.800 3.800  ;
    END
  END Y
  OBS
    VIA 1.800 22.500  dcont ;
    VIA 1.800 20.500  dcont ;
    VIA 1.800 3.800  dcont ;
    VIA 1.800 24.500  dcont ;
    VIA 4.800 22.500  dcont ;
    VIA 4.800 20.500  dcont ;
    VIA 4.800 24.500  dcont ;
    VIA 7.800 24.500  dcont ;
    VIA 7.800 22.500  dcont ;
    VIA 7.800 20.500  dcont ;
    VIA 8.800 3.800  dcont ;
    VIA 10.800 24.500  dcont ;
    VIA 10.800 22.500  dcont ;
    VIA 10.800 20.500  dcont ;
    VIA 11.800 3.800  dcont ;
    VIA 13.800 20.500  dcont ;
    VIA 13.800 22.500  dcont ;
    VIA 13.800 24.500  dcont ;
    VIA 5.000 13.500  pcont ;
    VIA 5.500 29.500  nsubcont ;
    VIA 8.000 10.700  pcont ;
    VIA 11.300 10.500  pcont ;
    VIA 2.000 10.700  pcont ;
    VIA 5.000 0.500  psubcont ;
    VIA 2.000 10.700  Via ;
    VIA 8.000 10.700  Via ;
    VIA 5.000 13.500  Via ;
    VIA 14.000 13.700  Via ;
  END
END an31

MACRO dcont
  CLASS BLOCK ;
END dcont

MACRO pcont
  CLASS BLOCK ;
END pcont

MACRO nsubcont
  CLASS BLOCK ;
  OBS
    VIA 0.000 0.000  dcont ;
  END
END nsubcont

MACRO psubcont
  CLASS BLOCK ;
  OBS
    VIA 0.000 0.000  dcont ;
  END
END psubcont

MACRO Via
  CLASS BLOCK ;
END Via


END LIBRARY
