VERSION 5.3 ;

NAMESCASESENSITIVE ON ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS











MACRO na222LEF
  CLASS BLOCK ;
  PIN A0
    DIRECTION INPUT ;
    PORT
      LAYER POL ;
        POLYGON 1.000 16.500  1.000 14.500  2.000 14.500  2.000 7.800  2.800 
        7.800  2.800 3.500  3.800 3.500  3.800 8.800  3.000 8.800  3.000 
        17.100  4.800 17.100  4.800 28.600  3.800 28.600  3.800 18.100  2.000 
        18.100  2.000 16.500  1.000 16.500  ;
    END
    PORT
      LAYER ML1 ;
        POLYGON 1.000 14.500  1.000 16.500  3.000 16.500  3.000 14.500  1.000 
        14.500  ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER POL ;
        POLYGON 4.000 12.300  4.000 10.300  5.000 10.300  5.000 9.500  5.800 
        9.500  5.800 3.500  6.800 3.500  6.800 10.500  6.000 10.500  6.000 
        15.000  6.800 15.000  6.800 26.500  5.800 26.500  5.800 16.000  5.000 
        16.000  5.000 12.300  4.000 12.300  ;
    END
    PORT
      LAYER ML1 ;
        POLYGON 4.000 10.300  4.000 12.300  6.000 12.300  6.000 10.300  4.000 
        10.300  ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    PORT
      LAYER POL ;
        POLYGON 10.000 16.500  10.000 14.500  11.800 14.500  11.800 3.500  
        12.800 3.500  12.800 16.200  12.000 16.200  12.000 16.500  11.800 
        16.500  11.800 26.500  10.800 26.500  10.800 16.500  10.000 16.500  ;
    END
    PORT
      LAYER ML1 ;
        POLYGON 10.000 14.500  10.000 16.500  12.000 16.500  12.000 14.500  
        10.000 14.500  ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER POL ;
        POLYGON 7.000 13.500  7.000 11.500  8.800 11.500  8.800 3.500  9.800 
        3.500  9.800 12.900  9.000 12.900  9.000 17.500  9.800 17.500  9.800 
        26.500  8.800 26.500  8.800 18.500  8.000 18.500  8.000 13.500  7.000 
        13.500  ;
    END
    PORT
      LAYER ML1 ;
        POLYGON 7.000 11.500  7.000 13.500  9.000 13.500  9.000 11.500  7.000 
        11.500  ;
    END
  END B1
  PIN VDD
    DIRECTION INOUT ;
    PORT
      LAYER ML1 ;
        POLYGON -0.500 30.500  -0.500 28.500  2.100 28.500  2.100 20.600  
        3.500 20.600  3.500 28.500  12.100 28.500  12.100 20.600  13.500 
        20.600  13.500 28.500  16.000 28.500  16.000 30.500  -0.500 30.500  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    PORT
      LAYER ML1 ;
        POLYGON -0.500 1.500  -0.500 -0.500  16.000 -0.500  16.000 1.500  
        5.300 1.500  5.300 6.000  4.300 6.000  4.300 1.500  -0.500 1.500  ;
    END
  END VSS
  PIN YB
    DIRECTION OUTPUT ;
    PORT
      LAYER ML1 ;
        POLYGON 10.300 8.500  10.300 5.000  11.300 5.000  11.300 7.500  14.000 
        7.500  14.000 10.500  15.000 10.500  15.000 12.500  14.000 12.500  
        14.000 18.500  8.300 18.500  8.300 20.600  8.500 20.600  8.500 25.200  
        7.100 25.200  7.100 20.600  7.300 20.600  7.300 17.500  13.000 17.500  
        13.000 8.500  10.300 8.500  ;
    END
  END YB
  OBS
    LAYER CNT ;
      POLYGON 10.300 5.000  10.300 6.000  11.300 6.000  11.300 5.000  10.300 
      5.000  ;
      POLYGON 12.300 20.000  12.300 21.000  13.300 21.000  13.300 20.000  
      12.300 20.000  ;
      POLYGON 12.300 22.000  12.300 23.000  13.300 23.000  13.300 22.000  
      12.300 22.000  ;
      POLYGON 12.300 24.000  12.300 25.000  13.300 25.000  13.300 24.000  
      12.300 24.000  ;
      POLYGON 13.300 5.000  13.300 6.000  14.300 6.000  14.300 5.000  13.300 
      5.000  ;
      POLYGON 10.500 15.000  10.500 16.000  11.500 16.000  11.500 15.000  
      10.500 15.000  ;
      POLYGON 7.500 12.000  7.500 13.000  8.500 13.000  8.500 12.000  7.500 
      12.000  ;
      POLYGON 9.700 29.000  9.700 30.000  10.700 30.000  10.700 29.000  9.700 
      29.000  ;
      POLYGON 4.500 10.800  4.500 11.800  5.500 11.800  5.500 10.800  4.500 
      10.800  ;
      POLYGON 1.500 15.000  1.500 16.000  2.500 16.000  2.500 15.000  1.500 
      15.000  ;
      POLYGON 9.700 0.000  9.700 1.000  10.700 1.000  10.700 0.000  9.700 
      0.000  ;
      POLYGON 7.300 5.000  7.300 6.000  8.300 6.000  8.300 5.000  7.300 5.000  ;
      
      POLYGON 7.300 20.000  7.300 21.000  8.300 21.000  8.300 20.000  7.300 
      20.000  ;
      POLYGON 7.300 22.000  7.300 23.000  8.300 23.000  8.300 22.000  7.300 
      22.000  ;
      POLYGON 7.300 24.000  7.300 25.000  8.300 25.000  8.300 24.000  7.300 
      24.000  ;
      POLYGON 4.300 5.000  4.300 6.000  5.300 6.000  5.300 5.000  4.300 5.000  ;
      
      POLYGON 2.300 24.000  2.300 25.000  3.300 25.000  3.300 24.000  2.300 
      24.000  ;
      POLYGON 2.300 20.000  2.300 21.000  3.300 21.000  3.300 20.000  2.300 
      20.000  ;
      POLYGON 2.300 22.000  2.300 23.000  3.300 23.000  3.300 22.000  2.300 
      22.000  ;
      POLYGON 1.300 5.000  1.300 6.000  2.300 6.000  2.300 5.000  1.300 5.000  ;
      
    LAYER FRAME ;
      RECT -0.500 28.500  16.000 30.500  ;
      RECT -0.500 -0.500  16.000 1.500  ;
      POLYGON 0.000 0.000  15.500 0.000  15.500 30.000  0.000 30.000  0.000 
      0.000  ;
    LAYER ML1 ;
      POLYGON 4.000 10.300  4.000 12.300  6.000 12.300  6.000 10.300  4.000 
      10.300  ;
      POLYGON 1.000 14.500  1.000 16.500  3.000 16.500  3.000 14.500  1.000 
      14.500  ;
      RECT 9.200 -0.500  11.200 1.500  ;
      POLYGON 7.000 11.500  7.000 13.500  9.000 13.500  9.000 11.500  7.000 
      11.500  ;
      POLYGON 10.000 14.500  10.000 16.500  12.000 16.500  12.000 14.500  
      10.000 14.500  ;
      RECT 1.000 14.500  3.000 16.500  ;
      RECT 4.000 10.300  6.000 12.300  ;
      RECT 9.200 28.500  11.200 30.500  ;
      RECT 7.000 11.500  9.000 13.500  ;
      RECT 10.000 14.500  12.000 16.500  ;
      RECT 12.800 4.500  14.800 6.500  ;
      RECT 11.800 23.500  13.800 25.500  ;
      RECT 11.800 21.500  13.800 23.500  ;
      RECT 11.800 19.500  13.800 21.500  ;
      RECT 9.800 4.500  11.800 6.500  ;
      RECT 6.800 4.500  8.800 6.500  ;
      RECT 6.800 19.500  8.800 21.500  ;
      RECT 6.800 21.500  8.800 23.500  ;
      RECT 6.800 23.500  8.800 25.500  ;
      RECT 3.800 4.500  5.800 6.500  ;
      RECT 1.800 23.500  3.800 25.500  ;
      RECT 1.800 19.500  3.800 21.500  ;
      RECT 1.800 21.500  3.800 23.500  ;
      RECT 0.800 4.500  2.800 6.500  ;
      POLYGON -0.500 30.500  -0.500 28.500  2.100 28.500  2.100 20.600  3.500 
      20.600  3.500 28.500  12.100 28.500  12.100 20.600  13.500 20.600  
      13.500 28.500  16.000 28.500  16.000 30.500  -0.500 30.500  ;
      POLYGON -0.500 1.500  -0.500 -0.500  16.000 -0.500  16.000 1.500  5.300 
      1.500  5.300 6.000  4.300 6.000  4.300 1.500  -0.500 1.500  ;
      POLYGON 1.300 8.500  1.300 5.000  2.300 5.000  2.300 7.500  7.300 7.500  
      7.300 2.500  14.300 2.500  14.300 6.000  13.300 6.000  13.300 3.500  
      8.300 3.500  8.300 8.500  1.300 8.500  ;
      POLYGON 10.300 8.500  10.300 5.000  11.300 5.000  11.300 7.500  14.000 
      7.500  14.000 10.500  15.000 10.500  15.000 12.500  14.000 12.500  
      14.000 18.500  8.300 18.500  8.300 20.600  8.500 20.600  8.500 25.200  
      7.100 25.200  7.100 20.600  7.300 20.600  7.300 17.500  13.000 17.500  
      13.000 8.500  10.300 8.500  ;
    LAYER ML2 ;
      POLYGON 13.000 12.500  13.000 10.500  15.000 10.500  15.000 12.500  
      13.000 12.500  ;
      POLYGON 10.000 14.500  10.000 16.500  12.000 16.500  12.000 14.500  
      10.000 14.500  ;
      POLYGON 7.000 11.500  7.000 13.500  9.000 13.500  9.000 11.500  7.000 
      11.500  ;
      POLYGON 4.000 10.300  4.000 12.300  6.000 12.300  6.000 10.300  4.000 
      10.300  ;
      POLYGON 1.000 14.500  1.000 16.500  3.000 16.500  3.000 14.500  1.000 
      14.500  ;
    LAYER POL ;
      POLYGON 10.000 16.500  10.000 14.500  11.800 14.500  11.800 3.500  
      12.800 3.500  12.800 16.200  12.000 16.200  12.000 16.500  11.800 16.500 
       11.800 26.500  10.800 26.500  10.800 16.500  10.000 16.500  ;
      POLYGON 7.000 13.500  7.000 11.500  8.800 11.500  8.800 3.500  9.800 
      3.500  9.800 12.900  9.000 12.900  9.000 17.500  9.800 17.500  9.800 
      26.500  8.800 26.500  8.800 18.500  8.000 18.500  8.000 13.500  7.000 
      13.500  ;
      POLYGON 4.000 12.300  4.000 10.300  5.000 10.300  5.000 9.500  5.800 
      9.500  5.800 3.500  6.800 3.500  6.800 10.500  6.000 10.500  6.000 
      15.000  6.800 15.000  6.800 26.500  5.800 26.500  5.800 16.000  5.000 
      16.000  5.000 12.300  4.000 12.300  ;
      POLYGON 1.000 16.500  1.000 14.500  2.000 14.500  2.000 7.800  2.800 
      7.800  2.800 3.500  3.800 3.500  3.800 8.800  3.000 8.800  3.000 17.100  
      4.800 17.100  4.800 28.600  3.800 28.600  3.800 18.100  2.000 18.100  
      2.000 16.500  1.000 16.500  ;
    LAYER VIA1 ;
      POLYGON 10.500 15.000  10.500 16.000  11.500 16.000  11.500 15.000  
      10.500 15.000  ;
      POLYGON 7.500 12.000  7.500 13.000  8.500 13.000  8.500 12.000  7.500 
      12.000  ;
      POLYGON 4.500 10.800  4.500 11.800  5.500 11.800  5.500 10.800  4.500 
      10.800  ;
      POLYGON 13.500 11.000  13.500 12.000  14.500 12.000  14.500 11.000  
      13.500 11.000  ;
      POLYGON 1.500 15.000  1.500 16.000  2.500 16.000  2.500 15.000  1.500 
      15.000  ;
  END
END na222LEF


END LIBRARY
