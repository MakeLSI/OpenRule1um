VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO dff1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 52.000 BY 30.000 ;
  SYMMETRY X Y ;
  SITE unit ;
  
  PIN CK
    USE SIGNAL ; ;
    PORT
      LAYER ML2 ;
        POLYGON 3.300 9.000  3.300 11.000  5.300 11.000  5.300 9.000  3.300 
        9.000  ;
    END
    PORT
      LAYER ML1 ;
        POLYGON 3.300 9.000  3.300 11.000  5.300 11.000  5.300 9.000  3.300 
        9.000  ;
    END
  END CK
  PIN D
    USE SIGNAL ; ;
    PORT
      LAYER ML1 ;
        POLYGON 11.000 9.000  11.000 11.000  13.000 11.000  13.000 9.000  
        11.000 9.000  ;
    END
    PORT
      LAYER ML2 ;
        POLYGON 11.000 9.000  11.000 11.000  13.000 11.000  13.000 9.000  
        11.000 9.000  ;
    END
  END D
  PIN Q
    USE SIGNAL ; ;
    PORT
      LAYER ML1 ;
        WIDTH 1.000  ;
        PATH 50.800 3.300 50.800 26.000  ;
    END
    PORT
      LAYER ML1 ;
        POLYGON 49.500 10.500  49.500 12.500  51.500 12.500  51.500 10.500  
        49.500 10.500  ;
    END
    PORT
      LAYER ML2 ;
        POLYGON 49.500 10.500  49.500 12.500  51.500 12.500  51.500 10.500  
        49.500 10.500  ;
    END
  END Q
  PIN VDD
    USE POWER ;
    PORT
      LAYER ML1 ;
        RECT -0.500 28.500  52.500 30.500  ;
    END
  END VDD
  PIN VSS
     USE GROUND ;
    PORT
      LAYER ML1 ;
        RECT -0.500 -0.500  52.500 1.500  ;
    END
  END VSS
  OBS

    LAYER ML1 ;
      WIDTH 1.400  ;
      PATH 1.800 22.600 1.800 25.800  ;

      WIDTH 1.400  ;
      PATH 50.300 22.600 50.300 25.800  ;
      WIDTH 1.000  ;
      PATH 1.800 3.800 1.800 21.800  ;
      WIDTH 1.000  ;
      PATH 5.800 18.800 1.800 18.800  ;
      WIDTH 1.000  ;
      PATH 5.300 13.000 1.800 13.000  ;
      WIDTH 1.000  ;
      PATH 5.800 6.800 1.800 6.800  ;
      WIDTH 1.000  ;
      PATH 8.300 25.800 8.300 16.200  ;
      WIDTH 1.000  ;
      PATH 14.800 6.800 8.300 6.800  ;
      WIDTH 1.000  ;
      PATH 8.300 3.600 8.300 9.500 7.800 9.500 7.800 16.200 31.300 16.200  ;
      WIDTH 1.000  ;
      PATH 16.300 21.800 16.300 18.800 22.300 18.800  ;
      WIDTH 1.000  ;
      PATH 26.800 19.200 25.000 19.200 25.000 21.300 24.300 21.300 24.300 
      21.800  ;
      WIDTH 1.000  ;
      PATH 38.800 19.200 32.800 19.200 32.800 21.800  ;
      WIDTH 1.000  ;
      PATH 41.300 25.800 41.300 3.700  ;
      WIDTH 1.000  ;
      PATH 45.300 8.800 41.300 8.800  ;
      WIDTH 1.000  ;
      PATH 36.800 14.000 41.300 14.000  ;
      WIDTH 1.000  ;
      PATH 45.300 17.200 41.300 17.200  ;
      WIDTH 1.000  ;
      PATH 20.300 6.800 26.800 6.800  ;
      WIDTH 1.000  ;
      PATH 24.300 6.800 24.300 3.700  ;
      WIDTH 1.000  ;
      PATH 32.800 3.800 32.800 6.800 38.800 6.800  ;
      WIDTH 1.000  ;
      PATH 44.300 3.800 44.300 6.300 48.000 6.300 48.000 19.400 44.200 19.400 
      44.200 21.800  ;
      WIDTH 1.000  ;
      PATH 50.800 3.300 50.800 26.000  ;
      WIDTH 1.400  ;
      PATH 7.800 22.600 7.800 25.800  ;
      WIDTH 1.400  ;
      PATH 16.300 22.600 16.300 25.800  ;
      WIDTH 1.400  ;
      PATH 24.300 22.600 24.300 25.800  ;
      WIDTH 1.400  ;
      PATH 32.800 22.600 32.800 25.800  ;
      WIDTH 1.400  ;
      PATH 40.800 22.600 40.800 25.800  ;
      WIDTH 1.400  ;
      PATH 44.300 22.600 44.300 25.800  ;
      WIDTH 1.400  ;
      PATH 50.300 22.600 50.300 25.800  ;

      WIDTH 1.400  ;
      PATH 4.800 3.800 4.800 1.500  ;
      WIDTH 1.400  ;
      PATH 11.300 3.800 11.300 1.500  ;
      WIDTH 1.400  ;
      PATH 21.300 3.800 21.300 1.500  ;
      WIDTH 1.400  ;
      PATH 27.800 3.800 27.800 1.500  ;
      WIDTH 1.400  ;
      PATH 37.800 3.800 37.800 1.500  ;
      WIDTH 1.400  ;
      PATH 47.300 3.800 47.300 1.500  ;
      WIDTH 1.400  ;
      PATH 4.800 21.800 4.800 28.500  ;
      WIDTH 1.400  ;
      PATH 11.300 21.800 11.300 28.500  ;
      WIDTH 1.400  ;
      PATH 21.300 21.800 21.300 28.500  ;
      WIDTH 1.400  ;
      PATH 27.800 21.800 27.800 28.500  ;
      WIDTH 1.400  ;
      PATH 37.800 21.800 37.800 28.500  ;
      WIDTH 1.400  ;
      PATH 47.300 21.800 47.300 28.500  ;

      WIDTH 1.000  ;
      PATH 10.300 13.000 34.000 13.000  ;
      WIDTH 1.000  ;
      PATH 22.300 10.000 16.800 10.000 16.800 4.300  ;

    VIA 22.300 18.700  pcont ;
    VIA 20.300 6.800  pcont ;
    VIA 17.300 16.000  pcont ;
    VIA 15.300 13.000  pcont ;
    VIA 14.800 6.800  pcont ;
    VIA 5.800 18.800  pcont ;
    VIA 10.300 13.000  pcont ;
    VIA 5.300 13.000  pcont ;
    VIA 5.800 6.800  pcont ;
    VIA 4.300 10.000  pcont ;
    VIA 12.000 10.000  pcont ;
    VIA 22.300 10.000  pcont ;
    VIA 26.800 6.800  pcont ;
    VIA 26.800 18.700  pcont ;
    VIA 28.800 13.000  pcont ;
    VIA 31.800 16.700  pcont ;
    VIA 33.800 13.700  pcont ;
    VIA 36.800 14.000  pcont ;
    VIA 38.800 6.800  pcont ;
    VIA 38.800 18.700  pcont ;
    VIA 45.300 8.800  pcont ;
    VIA 48.300 6.800  pcont ;
    VIA 48.300 18.900  pcont ;
    VIA 45.300 17.200  pcont ;
    VIA 46.000 0.500  psubcont ;
    VIA 27.700 0.500  psubcont ;
    VIA 10.200 0.500  psubcont ;
    VIA 27.700 29.500  nsubcont ;
    VIA 10.200 29.500  nsubcont ;
    VIA 46.000 29.500  nsubcont ;
    VIA 11.300 3.800  dcont ;
    VIA 16.300 3.800  dcont ;
    VIA 21.300 3.800  dcont ;
    VIA 24.300 3.800  dcont ;
    VIA 27.800 3.800  dcont ;
    VIA 32.800 3.800  dcont ;
    VIA 37.800 3.800  dcont ;
    VIA 40.800 3.800  dcont ;
    VIA 44.300 3.800  dcont ;
    VIA 47.300 3.800  dcont ;
    VIA 50.300 3.800  dcont ;
    VIA 7.800 3.800  dcont ;
    VIA 4.800 3.800  dcont ;
    VIA 1.800 3.800  dcont ;
    VIA 1.800 25.800  dcont ;
    VIA 1.800 23.800  dcont ;
    VIA 1.800 21.800  dcont ;
    VIA 4.800 21.800  dcont ;
    VIA 4.800 23.800  dcont ;
    VIA 4.800 25.800  dcont ;
    VIA 7.800 25.800  dcont ;
    VIA 7.800 23.800  dcont ;
    VIA 7.800 21.800  dcont ;
    VIA 11.300 21.800  dcont ;
    VIA 11.300 23.800  dcont ;
    VIA 11.300 25.800  dcont ;
    VIA 16.300 25.800  dcont ;
    VIA 16.300 23.800  dcont ;
    VIA 16.300 21.800  dcont ;
    VIA 21.300 21.800  dcont ;
    VIA 21.300 23.800  dcont ;
    VIA 21.300 25.800  dcont ;
    VIA 24.300 25.800  dcont ;
    VIA 24.300 23.800  dcont ;
    VIA 24.300 21.800  dcont ;
    VIA 27.800 21.800  dcont ;
    VIA 27.800 23.800  dcont ;
    VIA 27.800 25.800  dcont ;
    VIA 32.800 25.800  dcont ;
    VIA 32.800 23.800  dcont ;
    VIA 32.800 21.800  dcont ;
    VIA 37.800 21.800  dcont ;
    VIA 37.800 23.800  dcont ;
    VIA 37.800 25.800  dcont ;
    VIA 40.800 25.800  dcont ;
    VIA 40.800 23.800  dcont ;
    VIA 40.800 21.800  dcont ;
    VIA 44.300 25.800  dcont ;
    VIA 44.300 23.800  dcont ;
    VIA 44.300 21.800  dcont ;
    VIA 47.300 21.800  dcont ;
    VIA 47.300 23.800  dcont ;
    VIA 47.300 25.800  dcont ;
    VIA 50.300 25.800  dcont ;
    VIA 50.300 23.800  dcont ;
    VIA 50.300 21.800  dcont ;
  END
END dff1

MACRO pcont
  CLASS CORE ;
  OBS
    LAYER ML1 ;
      RECT -1.000 -1.000  1.000 1.000  ;
  END
END pcont

MACRO psubcont
  CLASS CORE ;
  OBS
    LAYER ML1 ;
      RECT -1.000 -1.000  1.000 1.000  ;
  END
END psubcont

MACRO nsubcont
  CLASS CORE ;
  OBS
    LAYER ML1 ;
      RECT -1.000 -1.000  1.000 1.000  ;
  END
END nsubcont

MACRO dcont
  CLASS CORE ;
  OBS
    LAYER ML1 ;
      RECT -1.000 -1.000  1.000 1.000  ;
  END
END dcont


END LIBRARY
