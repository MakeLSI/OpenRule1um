VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO na222
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 15.500 BY 30.000 ;
  SYMMETRY X Y ;
  SITE unit ;
 
  PIN A0
    USE SIGNAL ;
    PORT
      LAYER ML2 ;
        POLYGON 1.000 14.500  1.000 16.500  3.000 16.500  3.000 14.500  1.000 
        14.500  ;
    END
    PORT
      LAYER ML1 ;
        POLYGON 1.000 14.500  1.000 16.500  3.000 16.500  3.000 14.500  1.000 
        14.500  ;
    END
  END A0
  PIN A1
    USE SIGNAL ;
    PORT
      LAYER ML2 ;
        POLYGON 4.000 10.300  4.000 12.300  6.000 12.300  6.000 10.300  4.000 
        10.300  ;
    END
    PORT
      LAYER ML1 ;
        POLYGON 4.000 10.300  4.000 12.300  6.000 12.300  6.000 10.300  4.000 
        10.300  ;
    END
  END A1
  PIN B0
    USE SIGNAL ;
    PORT
      LAYER ML2 ;
        POLYGON 10.000 14.500  10.000 16.500  12.000 16.500  12.000 14.500  
        10.000 14.500  ;
    END
    PORT
      LAYER ML1 ;
        POLYGON 10.000 14.500  10.000 16.500  12.000 16.500  12.000 14.500  
        10.000 14.500  ;
    END
  END B0
  PIN B1
    USE SIGNAL ;
    PORT
      LAYER ML2 ;
        POLYGON 7.000 11.500  7.000 13.500  9.000 13.500  9.000 11.500  7.000 
        11.500  ;
    END
    PORT
      LAYER ML1 ;
        POLYGON 7.000 11.500  7.000 13.500  9.000 13.500  9.000 11.500  7.000 
        11.500  ;
    END
  END B1
  PIN VDD
    USE POWER ;
    PORT
      LAYER ML1 ;
        RECT -0.500 28.500  16.000 30.500  ;
    END
  END VDD
  PIN VSS
     USE GROUND ;
    PORT
      LAYER ML1 ;
        RECT -0.500 -0.500  16.000 1.500  ;
    END
  END VSS
  PIN YB
    USE SIGNAL ;
    PORT
      LAYER ML1 ;
        WIDTH 1.000  ;
        PATH 7.800 20.500 7.800 18.000 13.500 18.000 13.500 8.000 10.800 8.000 
        10.800 5.500  ;
    END
    PORT
      LAYER ML1 ;
        POLYGON 13.000 10.500  13.000 12.500  15.000 12.500  15.000 10.500  
        13.000 10.500  ;
    END
    PORT
      LAYER ML2 ;
        POLYGON 13.000 10.500  13.000 12.500  15.000 12.500  15.000 10.500  
        13.000 10.500  ;
    END
  END YB
  OBS

    LAYER ML1 ;
      POLYGON 4.000 10.300  4.000 12.300  6.000 12.300  6.000 10.300  4.000 
      10.300  ;
      POLYGON 1.000 14.500  1.000 16.500  3.000 16.500  3.000 14.500  1.000 
      14.500  ;
      POLYGON 13.000 10.500  13.000 12.500  15.000 12.500  15.000 10.500  
      13.000 10.500  ;
      WIDTH 1.000  ;
      PATH 13.800 5.500 13.800 3.000 7.800 3.000 7.800 8.000 1.800 8.000 1.800 
      5.500  ;
      WIDTH 1.000  ;
      PATH 4.800 1.000 4.800 5.500  ;
      WIDTH 1.400  ;
      PATH 2.800 21.300 2.800 28.500  ;

      WIDTH 1.000  ;
      PATH 7.800 20.500 7.800 18.000 13.500 18.000 13.500 8.000 10.800 8.000 
      10.800 5.500  ;
      WIDTH 1.400  ;
      PATH 12.800 21.300 12.800 28.500  ;
      WIDTH 1.400  ;
      PATH 7.800 21.300 7.800 24.500  ;

    VIA 1.800 5.500  dcont ;
    VIA 2.800 22.500  dcont ;
    VIA 2.800 20.500  dcont ;
    VIA 2.800 24.500  dcont ;
    VIA 4.800 5.500  dcont ;
    VIA 7.800 24.500  dcont ;
    VIA 7.800 22.500  dcont ;
    VIA 7.800 20.500  dcont ;
    VIA 7.800 5.500  dcont ;
    VIA 10.800 5.500  dcont ;
    VIA 12.800 20.500  dcont ;
    VIA 12.800 22.500  dcont ;
    VIA 12.800 24.500  dcont ;
    VIA 13.800 5.500  dcont ;
    VIA 11.000 15.500  pcont ;
    VIA 8.000 12.500  pcont ;
    VIA 10.200 29.500  nsubcont ;
    VIA 5.000 11.300  pcont ;
    VIA 2.000 15.500  pcont ;
    VIA 10.200 0.500  psubcont ;
  END
END na222

MACRO dcont
  CLASS CORE ;
  OBS
    LAYER ML1 ;
      RECT -1.000 -1.000  1.000 1.000  ;
  END
END dcont

MACRO pcont
  CLASS CORE ;
  OBS
    LAYER ML1 ;
      RECT -1.000 -1.000  1.000 1.000  ;
  END
END pcont

MACRO nsubcont
  CLASS CORE ;
  OBS
    LAYER ML1 ;
      RECT -1.000 -1.000  1.000 1.000  ;
  END
END nsubcont

MACRO psubcont
  CLASS CORE ;
  OBS
    LAYER ML1 ;
      RECT -1.000 -1.000  1.000 1.000  ;
  END
END psubcont


END LIBRARY
