VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO exor
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 21.000 BY 30.000 ;
  SYMMETRY X Y ;
  SITE unit ;
 
  PIN A
    USE SIGNAL ;
    PORT
      LAYER ML1 ;
        WIDTH 1.000  ;
        PATH 7.000 14.700 14.800 14.700  ;
    END
    PORT
      LAYER ML1 ;
        POLYGON 6.000 13.700  6.000 15.700  8.000 15.700  8.000 13.700  6.000 
        13.700  ;
    END
    PORT
      LAYER ML2 ;
        POLYGON 6.000 13.700  6.000 15.700  8.000 15.700  8.000 13.700  6.000 
        13.700  ;
    END
  END A
  PIN B
    USE SIGNAL ;
    PORT
      LAYER ML1 ;
        WIDTH 1.000  ;
        PATH 4.000 10.700 11.300 10.700  ;
    END
    PORT
      LAYER ML1 ;
        POLYGON 3.000 9.700  3.000 11.700  5.000 11.700  5.000 9.700  3.000 
        9.700  ;
    END
    PORT
      LAYER ML2 ;
        POLYGON 3.000 9.700  3.000 11.700  5.000 11.700  5.000 9.700  3.000 
        9.700  ;
    END
  END B
  PIN VDD
    USE POWER ;
    PORT
      LAYER ML1 ;
        RECT -0.500 28.500  21.500 30.500  ;
    END
  END VDD
  PIN VSS
    USE GROUND ;
    PORT
      LAYER ML1 ;
        RECT -0.500 -0.500  21.500 1.500  ;
    END
  END VSS
  PIN Y
    USE SIGNAL ;
    PORT
      LAYER ML1 ;
        WIDTH 1.000  ;
        PATH 19.300 21.800 19.300 5.700 15.300 5.700 15.300 3.800  ;
    END
    PORT
      LAYER ML2 ;
        POLYGON 18.500 12.700  18.500 14.700  20.500 14.700  20.500 12.700  
        18.500 12.700  ;
    END
    PORT
      LAYER ML1 ;
        POLYGON 18.500 12.700  18.500 14.700  20.500 14.700  20.500 12.700  
        18.500 12.700  ;
    END
  END Y
  OBS

    LAYER ML1 ;
      WIDTH 1.400  ;
      PATH 1.800 22.600 1.800 25.800  ;
      WIDTH 1.000  ;
      PATH 1.800 1.000 1.800 3.800  ;
      WIDTH 1.000  ;
      PATH 4.800 8.200 4.800 3.800  ;
      WIDTH 1.400  ;
      PATH 6.800 22.600 6.800 28.500  ;
      WIDTH 1.000  ;
      PATH 4.000 10.700 11.300 10.700  ;
      WIDTH 1.000  ;
      PATH 7.800 1.000 7.800 3.800  ;
      WIDTH 1.000  ;
      PATH 1.800 25.800 1.800 19.000 1.500 19.000 1.500 8.200 16.800 8.200  ;
      WIDTH 1.000  ;
      PATH 10.300 1.000 10.300 3.800  ;

      WIDTH 1.000  ;
      PATH 7.000 14.700 14.800 14.700  ;
      WIDTH 1.400  ;
      PATH 13.300 22.600 13.300 28.500  ;
      WIDTH 1.400  ;
      PATH 16.300 25.800 16.300 19.500 10.300 19.500 10.300 25.100  ;
      WIDTH 1.000  ;
      PATH 19.300 21.800 19.300 5.700 15.300 5.700 15.300 3.800  ;
      WIDTH 1.000  ;
      PATH 18.300 1.000 18.300 3.800  ;
      WIDTH 1.400  ;
      PATH 19.300 21.800 19.300 25.800  ;

    VIA 1.800 23.800  dcont ;
    VIA 1.800 21.800  dcont ;
    VIA 1.800 3.800  dcont ;
    VIA 1.800 25.800  dcont ;
    VIA 4.800 3.800  dcont ;
    VIA 6.800 23.800  dcont ;
    VIA 6.800 21.800  dcont ;
    VIA 6.800 25.800  dcont ;
    VIA 7.800 3.800  dcont ;
    VIA 10.300 21.800  dcont ;
    VIA 10.300 23.800  dcont ;
    VIA 10.300 25.800  dcont ;
    VIA 10.300 3.800  dcont ;
    VIA 13.300 21.800  dcont ;
    VIA 13.300 23.800  dcont ;
    VIA 13.300 25.800  dcont ;
    VIA 15.300 3.800  dcont ;
    VIA 16.300 21.800  dcont ;
    VIA 16.300 25.800  dcont ;
    VIA 16.300 23.800  dcont ;
    VIA 18.300 3.800  dcont ;
    VIA 19.300 23.800  dcont ;
    VIA 19.300 21.800  dcont ;
    VIA 19.300 25.800  dcont ;
    VIA 7.000 14.700  pcont ;
    VIA 10.200 29.500  nsubcont ;
    VIA 17.000 8.200  pcont ;
    VIA 14.300 14.700  pcont ;
    VIA 4.000 10.700  pcont ;
    VIA 11.300 10.700  pcont ;
    VIA 10.200 0.500  psubcont ;
  END
END exor

MACRO dcont
  CLASS CORE ;
  OBS
    LAYER ML1 ;
      RECT -1.000 -1.000  1.000 1.000  ;
  END
END dcont

MACRO pcont
  CLASS CORE ;
  OBS
    LAYER ML1 ;
      RECT -1.000 -1.000  1.000 1.000  ;
  END
END pcont

MACRO nsubcont
  CLASS CORE ;
  OBS
    LAYER ML1 ;
      RECT -1.000 -1.000  1.000 1.000  ;
  END
END nsubcont

MACRO psubcont
  CLASS CORE ;
  OBS
    LAYER ML1 ;
      RECT -1.000 -1.000  1.000 1.000  ;
  END
END psubcont


END LIBRARY
