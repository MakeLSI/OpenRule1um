VERSION 5.3 ;

NAMESCASESENSITIVE ON ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS











MACRO exnrLEF
  CLASS BLOCK ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER POL ;
        POLYGON 4.800 8.000  4.800 1.700  5.800 1.700  5.800 7.000  7.000 
        7.000  7.000 13.700  8.000 13.700  8.000 15.700  7.000 15.700  7.000 
        18.000  6.800 18.000  6.800 27.800  5.800 27.800  5.800 17.000  6.000 
        17.000  6.000 8.000  4.800 8.000  ;
    END
    PORT
      LAYER ML1 ;
        POLYGON 6.000 15.700  6.000 13.700  8.000 13.700  8.000 14.200  13.300 
        14.200  13.300 13.700  15.300 13.700  15.300 15.700  13.300 15.700  
        13.300 15.200  8.000 15.200  8.000 15.700  6.000 15.700  ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER POL ;
        POLYGON 2.800 27.800  2.800 1.700  3.800 1.700  3.800 10.700  5.000 
        10.700  5.000 12.700  3.800 12.700  3.800 27.800  2.800 27.800  ;
    END
    PORT
      LAYER ML1 ;
        POLYGON 3.000 12.700  3.000 10.700  5.000 10.700  5.000 11.200  10.300 
        11.200  10.300 10.700  12.300 10.700  12.300 12.700  10.300 12.700  
        10.300 12.200  5.000 12.200  5.000 12.700  3.000 12.700  ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    PORT
      LAYER ML1 ;
        POLYGON -0.500 30.500  -0.500 28.500  1.100 28.500  1.100 21.900  
        2.500 21.900  2.500 28.500  7.100 28.500  7.100 21.900  8.500 21.900  
        8.500 28.500  10.600 28.500  10.600 21.900  12.000 21.900  12.000 
        28.500  18.600 28.500  18.600 21.900  20.000 21.900  20.000 28.500  
        21.500 28.500  21.500 30.500  -0.500 30.500  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    PORT
      LAYER ML1 ;
        POLYGON -0.500 1.500  -0.500 -0.500  21.500 -0.500  21.500 1.500  
        13.800 1.500  13.800 4.200  12.800 4.200  12.800 1.500  7.300 1.500  
        7.300 4.200  6.300 4.200  6.300 1.500  -0.500 1.500  ;
    END
  END VSS
  PIN YB
    DIRECTION OUTPUT ;
    PORT
      LAYER ML1 ;
        POLYGON 18.800 6.700  18.800 3.200  19.800 3.200  19.800 5.700  20.300 
        5.700  20.300 12.500  20.500 12.500  20.500 14.500  20.300 14.500  
        20.300 18.000  16.800 18.000  16.800 21.100  17.000 21.100  17.000 
        26.500  15.600 26.500  15.600 21.100  15.800 21.100  15.800 17.000  
        19.300 17.000  19.300 14.500  18.500 14.500  18.500 12.500  19.300 
        12.500  19.300 6.700  18.800 6.700  ;
    END
  END YB
  OBS
    LAYER CNT ;
      POLYGON 18.800 23.300  18.800 24.300  19.800 24.300  19.800 23.300  
      18.800 23.300  ;
      POLYGON 18.800 21.300  18.800 22.300  19.800 22.300  19.800 21.300  
      18.800 21.300  ;
      POLYGON 18.800 25.300  18.800 26.300  19.800 26.300  19.800 25.300  
      18.800 25.300  ;
      POLYGON 18.800 3.200  18.800 4.200  19.800 4.200  19.800 3.200  18.800 
      3.200  ;
      POLYGON 13.800 14.200  13.800 15.200  14.800 15.200  14.800 14.200  
      13.800 14.200  ;
      POLYGON 16.800 8.200  16.800 9.200  17.800 9.200  17.800 8.200  16.800 
      8.200  ;
      POLYGON 9.700 29.000  9.700 30.000  10.700 30.000  10.700 29.000  9.700 
      29.000  ;
      POLYGON 6.500 14.200  6.500 15.200  7.500 15.200  7.500 14.200  6.500 
      14.200  ;
      POLYGON 10.800 11.200  10.800 12.200  11.800 12.200  11.800 11.200  
      10.800 11.200  ;
      POLYGON 3.500 11.200  3.500 12.200  4.500 12.200  4.500 11.200  3.500 
      11.200  ;
      POLYGON 9.700 0.000  9.700 1.000  10.700 1.000  10.700 0.000  9.700 
      0.000  ;
      POLYGON 15.800 3.200  15.800 4.200  16.800 4.200  16.800 3.200  15.800 
      3.200  ;
      POLYGON 15.800 23.300  15.800 24.300  16.800 24.300  16.800 23.300  
      15.800 23.300  ;
      POLYGON 15.800 25.300  15.800 26.300  16.800 26.300  16.800 25.300  
      15.800 25.300  ;
      POLYGON 15.800 21.300  15.800 22.300  16.800 22.300  16.800 21.300  
      15.800 21.300  ;
      POLYGON 12.800 3.200  12.800 4.200  13.800 4.200  13.800 3.200  12.800 
      3.200  ;
      POLYGON 10.800 25.300  10.800 26.300  11.800 26.300  11.800 25.300  
      10.800 25.300  ;
      POLYGON 10.800 23.300  10.800 24.300  11.800 24.300  11.800 23.300  
      10.800 23.300  ;
      POLYGON 10.800 21.300  10.800 22.300  11.800 22.300  11.800 21.300  
      10.800 21.300  ;
      POLYGON 9.800 3.200  9.800 4.200  10.800 4.200  10.800 3.200  9.800 
      3.200  ;
      POLYGON 7.300 25.300  7.300 26.300  8.300 26.300  8.300 25.300  7.300 
      25.300  ;
      POLYGON 7.300 21.300  7.300 22.300  8.300 22.300  8.300 21.300  7.300 
      21.300  ;
      POLYGON 7.300 23.300  7.300 24.300  8.300 24.300  8.300 23.300  7.300 
      23.300  ;
      POLYGON 6.300 3.200  6.300 4.200  7.300 4.200  7.300 3.200  6.300 3.200  ;
      
      POLYGON 4.300 21.300  4.300 22.300  5.300 22.300  5.300 21.300  4.300 
      21.300  ;
      POLYGON 4.300 23.300  4.300 24.300  5.300 24.300  5.300 23.300  4.300 
      23.300  ;
      POLYGON 4.300 25.300  4.300 26.300  5.300 26.300  5.300 25.300  4.300 
      25.300  ;
      POLYGON 1.300 25.300  1.300 26.300  2.300 26.300  2.300 25.300  1.300 
      25.300  ;
      POLYGON 1.300 3.200  1.300 4.200  2.300 4.200  2.300 3.200  1.300 3.200  ;
      
      POLYGON 1.300 21.300  1.300 22.300  2.300 22.300  2.300 21.300  1.300 
      21.300  ;
      POLYGON 1.300 23.300  1.300 24.300  2.300 24.300  2.300 23.300  1.300 
      23.300  ;
    LAYER FRAME ;
      POLYGON -0.500 1.500  -0.500 -0.500  21.500 -0.500  21.500 1.500  -0.500 
      1.500  ;
      POLYGON 0.000 0.000  21.000 0.000  21.000 30.000  0.000 30.000  0.000 
      0.000  ;
      RECT -0.500 28.500  21.500 30.500  ;
    LAYER ML1 ;
      RECT 0.800 24.800  2.800 26.800  ;
      RECT 0.800 2.700  2.800 4.700  ;
      RECT 0.800 20.800  2.800 22.800  ;
      RECT 0.800 22.800  2.800 24.800  ;
      RECT 3.800 20.800  5.800 22.800  ;
      RECT 3.800 22.800  5.800 24.800  ;
      RECT 3.800 24.800  5.800 26.800  ;
      RECT 5.800 2.700  7.800 4.700  ;
      RECT 6.800 24.800  8.800 26.800  ;
      RECT 6.800 20.800  8.800 22.800  ;
      RECT 6.800 22.800  8.800 24.800  ;
      RECT 9.200 -0.500  11.200 1.500  ;
      RECT 9.200 28.500  11.200 30.500  ;
      RECT 9.300 2.700  11.300 4.700  ;
      RECT 10.300 24.800  12.300 26.800  ;
      RECT 10.300 22.800  12.300 24.800  ;
      RECT 10.300 20.800  12.300 22.800  ;
      RECT 12.300 2.700  14.300 4.700  ;
      RECT 15.300 2.700  17.300 4.700  ;
      RECT 15.300 22.800  17.300 24.800  ;
      RECT 15.300 24.800  17.300 26.800  ;
      RECT 15.300 20.800  17.300 22.800  ;
      RECT 18.300 2.700  20.300 4.700  ;
      RECT 18.300 24.800  20.300 26.800  ;
      RECT 18.300 20.800  20.300 22.800  ;
      RECT 18.300 22.800  20.300 24.800  ;
      POLYGON -0.500 30.500  -0.500 28.500  1.100 28.500  1.100 21.900  2.500 
      21.900  2.500 28.500  7.100 28.500  7.100 21.900  8.500 21.900  8.500 
      28.500  10.600 28.500  10.600 21.900  12.000 21.900  12.000 28.500  
      18.600 28.500  18.600 21.900  20.000 21.900  20.000 28.500  21.500 
      28.500  21.500 30.500  -0.500 30.500  ;
      POLYGON -0.500 1.500  -0.500 -0.500  21.500 -0.500  21.500 1.500  13.800 
      1.500  13.800 4.200  12.800 4.200  12.800 1.500  7.300 1.500  7.300 
      4.200  6.300 4.200  6.300 1.500  -0.500 1.500  ;
      POLYGON 1.000 19.500  1.000 5.500  1.300 5.500  1.300 3.200  2.300 3.200 
       2.300 6.500  2.000 6.500  2.000 8.200  16.300 8.200  16.300 7.700  
      18.300 7.700  18.300 9.700  16.300 9.700  16.300 9.200  2.000 9.200  
      2.000 18.500  5.300 18.500  5.300 26.300  4.300 26.300  4.300 19.500  
      1.000 19.500  ;
      POLYGON 3.000 12.700  3.000 10.700  5.000 10.700  5.000 11.200  10.300 
      11.200  10.300 10.700  12.300 10.700  12.300 12.700  10.300 12.700  
      10.300 12.200  5.000 12.200  5.000 12.700  3.000 12.700  ;
      POLYGON 6.000 15.700  6.000 13.700  8.000 13.700  8.000 14.200  13.300 
      14.200  13.300 13.700  15.300 13.700  15.300 15.700  13.300 15.700  
      13.300 15.200  8.000 15.200  8.000 15.700  6.000 15.700  ;
      POLYGON 9.800 6.700  9.800 3.200  10.800 3.200  10.800 5.700  15.800 
      5.700  15.800 3.200  16.800 3.200  16.800 6.700  9.800 6.700  ;
      POLYGON 18.800 6.700  18.800 3.200  19.800 3.200  19.800 5.700  20.300 
      5.700  20.300 12.500  20.500 12.500  20.500 14.500  20.300 14.500  
      20.300 18.000  16.800 18.000  16.800 21.100  17.000 21.100  17.000 
      26.500  15.600 26.500  15.600 21.100  15.800 21.100  15.800 17.000  
      19.300 17.000  19.300 14.500  18.500 14.500  18.500 12.500  19.300 
      12.500  19.300 6.700  18.800 6.700  ;
    LAYER ML2 ;
      POLYGON 6.000 15.700  6.000 13.700  8.000 13.700  8.000 15.700  6.000 
      15.700  ;
      POLYGON 3.000 12.700  3.000 10.700  5.000 10.700  5.000 12.700  3.000 
      12.700  ;
      POLYGON 18.500 12.500  18.500 14.500  20.500 14.500  20.500 12.500  
      18.500 12.500  ;
    LAYER POL ;
      POLYGON 16.300 9.700  16.300 7.700  17.300 7.700  17.300 1.900  18.300 
      1.900  18.300 27.600  17.300 27.600  17.300 9.700  16.300 9.700  ;
      POLYGON 13.300 15.700  13.300 13.700  14.300 13.700  14.300 1.900  
      15.300 1.900  15.300 27.600  14.300 27.600  14.300 15.700  13.300 15.700 
       ;
      POLYGON 10.300 12.700  10.300 10.700  11.300 10.700  11.300 1.900  
      12.300 1.900  12.300 17.500  13.300 17.500  13.300 27.600  12.300 27.600 
       12.300 18.500  11.300 18.500  11.300 12.700  10.300 12.700  ;
      POLYGON 4.800 8.000  4.800 1.700  5.800 1.700  5.800 7.000  7.000 7.000  
      7.000 13.700  8.000 13.700  8.000 15.700  7.000 15.700  7.000 18.000  
      6.800 18.000  6.800 27.800  5.800 27.800  5.800 17.000  6.000 17.000  
      6.000 8.000  4.800 8.000  ;
      POLYGON 2.800 27.800  2.800 1.700  3.800 1.700  3.800 10.700  5.000 
      10.700  5.000 12.700  3.800 12.700  3.800 27.800  2.800 27.800  ;
    LAYER VIA1 ;
      POLYGON 3.500 11.200  3.500 12.200  4.500 12.200  4.500 11.200  3.500 
      11.200  ;
      POLYGON 19.000 13.000  19.000 14.000  20.000 14.000  20.000 13.000  
      19.000 13.000  ;
      POLYGON 6.500 14.200  6.500 15.200  7.500 15.200  7.500 14.200  6.500 
      14.200  ;
  END
END exnrLEF


END LIBRARY
