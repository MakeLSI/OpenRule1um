VERSION 5.3 ;

NAMESCASESENSITIVE ON ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS











MACRO an41LEF
  CLASS BLOCK ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER POL ;
        POLYGON 1.000 17.500  1.000 15.500  2.000 15.500  2.000 6.500  2.800 
        6.500  2.800 1.700  3.800 1.700  3.800 7.500  3.000 7.500  3.000 
        15.500  3.800 15.500  3.800 26.500  2.800 26.500  2.800 17.500  1.000 
        17.500  ;
    END
    PORT
      LAYER ML1 ;
        POLYGON 1.000 15.500  1.000 17.500  3.000 17.500  3.000 15.500  1.000 
        15.500  ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER POL ;
        POLYGON 4.000 14.500  4.000 12.500  4.800 12.500  4.800 1.700  5.800 
        1.700  5.800 12.500  6.000 12.500  6.000 13.500  6.800 13.500  6.800 
        26.500  5.800 26.500  5.800 14.500  4.000 14.500  ;
    END
    PORT
      LAYER ML1 ;
        POLYGON 4.000 14.500  4.000 12.500  6.000 12.500  6.000 14.500  4.000 
        14.500  ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER POL ;
        POLYGON 6.800 11.500  6.800 1.700  7.800 1.700  7.800 9.700  9.000 
        9.700  9.000 11.700  8.800 11.700  8.800 16.500  9.800 16.500  9.800 
        26.500  8.800 26.500  8.800 17.500  7.800 17.500  7.800 11.700  7.000 
        11.700  7.000 11.500  6.800 11.500  ;
    END
    PORT
      LAYER ML1 ;
        POLYGON 7.000 9.700  7.000 11.700  9.000 11.700  9.000 9.700  7.000 
        9.700  ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER POL ;
        POLYGON 8.800 8.700  8.800 1.700  9.800 1.700  9.800 7.700  11.300 
        7.700  11.300 12.500  12.000 12.500  12.000 13.000  12.800 13.000  
        12.800 26.500  11.800 26.500  11.800 14.500  10.000 14.500  10.000 
        12.500  10.300 12.500  10.300 8.700  8.800 8.700  ;
    END
    PORT
      LAYER ML1 ;
        RECT 10.000 12.500  12.000 14.500  ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    PORT
      LAYER ML1 ;
        POLYGON -0.500 1.500  -0.500 -0.500  19.000 -0.500  19.000 1.500  
        2.300 1.500  2.300 4.200  1.300 4.200  1.300 1.500  -0.500 1.500  ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    PORT
      LAYER ML1 ;
        POLYGON 13.300 8.500  13.300 3.200  14.300 3.200  14.300 7.500  17.300 
        7.500  17.300 12.700  18.000 12.700  18.000 14.700  17.300 14.700  
        17.300 20.600  17.500 20.600  17.500 25.200  16.100 25.200  16.100 
        20.600  16.300 20.600  16.300 14.700  16.000 14.700  16.000 12.700  
        16.300 12.700  16.300 8.500  13.300 8.500  ;
    END
  END Y
  OBS
    LAYER CNT ;
      POLYGON 13.300 3.200  13.300 4.200  14.300 4.200  14.300 3.200  13.300 
      3.200  ;
      POLYGON 16.300 20.000  16.300 21.000  17.300 21.000  17.300 20.000  
      16.300 20.000  ;
      POLYGON 16.300 22.000  16.300 23.000  17.300 23.000  17.300 22.000  
      16.300 22.000  ;
      POLYGON 16.300 24.000  16.300 25.000  17.300 25.000  17.300 24.000  
      16.300 24.000  ;
      POLYGON 13.800 10.000  13.800 11.000  14.800 11.000  14.800 10.000  
      13.800 10.000  ;
      POLYGON 10.500 13.000  10.500 14.000  11.500 14.000  11.500 13.000  
      10.500 13.000  ;
      POLYGON 7.500 10.200  7.500 11.200  8.500 11.200  8.500 10.200  7.500 
      10.200  ;
      POLYGON 5.000 29.000  5.000 30.000  6.000 30.000  6.000 29.000  5.000 
      29.000  ;
      POLYGON 4.500 13.000  4.500 14.000  5.500 14.000  5.500 13.000  4.500 
      13.000  ;
      POLYGON 1.500 16.000  1.500 17.000  2.500 17.000  2.500 16.000  1.500 
      16.000  ;
      POLYGON 4.500 0.000  4.500 1.000  5.500 1.000  5.500 0.000  4.500 0.000  ;
      
      POLYGON 13.300 20.000  13.300 21.000  14.300 21.000  14.300 20.000  
      13.300 20.000  ;
      POLYGON 13.300 22.000  13.300 23.000  14.300 23.000  14.300 22.000  
      13.300 22.000  ;
      POLYGON 13.300 24.000  13.300 25.000  14.300 25.000  14.300 24.000  
      13.300 24.000  ;
      POLYGON 10.300 24.000  10.300 25.000  11.300 25.000  11.300 24.000  
      10.300 24.000  ;
      POLYGON 10.300 22.000  10.300 23.000  11.300 23.000  11.300 22.000  
      10.300 22.000  ;
      POLYGON 10.300 20.000  10.300 21.000  11.300 21.000  11.300 20.000  
      10.300 20.000  ;
      POLYGON 10.300 3.200  10.300 4.200  11.300 4.200  11.300 3.200  10.300 
      3.200  ;
      POLYGON 7.300 20.000  7.300 21.000  8.300 21.000  8.300 20.000  7.300 
      20.000  ;
      POLYGON 7.300 22.000  7.300 23.000  8.300 23.000  8.300 22.000  7.300 
      22.000  ;
      POLYGON 7.300 24.000  7.300 25.000  8.300 25.000  8.300 24.000  7.300 
      24.000  ;
      POLYGON 4.300 24.000  4.300 25.000  5.300 25.000  5.300 24.000  4.300 
      24.000  ;
      POLYGON 4.300 20.000  4.300 21.000  5.300 21.000  5.300 20.000  4.300 
      20.000  ;
      POLYGON 4.300 22.000  4.300 23.000  5.300 23.000  5.300 22.000  4.300 
      22.000  ;
      POLYGON 1.300 24.000  1.300 25.000  2.300 25.000  2.300 24.000  1.300 
      24.000  ;
      POLYGON 1.300 3.200  1.300 4.200  2.300 4.200  2.300 3.200  1.300 3.200  ;
      
      POLYGON 1.300 20.000  1.300 21.000  2.300 21.000  2.300 20.000  1.300 
      20.000  ;
      POLYGON 1.300 22.000  1.300 23.000  2.300 23.000  2.300 22.000  1.300 
      22.000  ;
    LAYER FRAME ;
      RECT -0.500 28.500  19.000 30.500  ;
      RECT -0.500 -0.500  19.000 1.500  ;
      POLYGON 0.000 0.000  18.500 0.000  18.500 30.000  0.000 30.000  0.000 
      0.000  ;
    LAYER ML1 ;
      RECT 0.800 23.500  2.800 25.500  ;
      RECT 0.800 2.700  2.800 4.700  ;
      RECT 0.800 19.500  2.800 21.500  ;
      RECT 0.800 21.500  2.800 23.500  ;
      POLYGON 1.000 15.500  1.000 17.500  3.000 17.500  3.000 15.500  1.000 
      15.500  ;
      RECT 1.000 15.500  3.000 17.500  ;
      RECT 3.800 23.500  5.800 25.500  ;
      RECT 3.800 19.500  5.800 21.500  ;
      RECT 3.800 21.500  5.800 23.500  ;
      RECT 4.000 -0.500  6.000 1.500  ;
      POLYGON 4.000 14.500  4.000 12.500  6.000 12.500  6.000 14.500  4.000 
      14.500  ;
      RECT 4.500 28.500  6.500 30.500  ;
      RECT 6.800 19.500  8.800 21.500  ;
      RECT 6.800 21.500  8.800 23.500  ;
      RECT 6.800 23.500  8.800 25.500  ;
      POLYGON 7.000 9.700  7.000 11.700  9.000 11.700  9.000 9.700  7.000 
      9.700  ;
      RECT 7.000 9.700  9.000 11.700  ;
      POLYGON -0.500 1.500  -0.500 -0.500  19.000 -0.500  19.000 1.500  2.300 
      1.500  2.300 4.200  1.300 4.200  1.300 1.500  -0.500 1.500  ;
      POLYGON -0.500 30.500  -0.500 28.500  1.100 28.500  1.100 20.600  2.500 
      20.600  2.500 28.500  7.100 28.500  7.100 20.600  8.500 20.600  8.500 
      28.500  13.100 28.500  13.100 20.600  14.500 20.600  14.500 28.500  
      19.000 28.500  19.000 30.500  -0.500 30.500  ;
      POLYGON 10.300 10.500  10.300 3.200  11.300 3.200  11.300 9.500  15.300 
      9.500  15.300 11.500  14.300 11.500  14.300 18.500  11.300 18.500  
      11.300 20.600  11.500 20.600  11.500 25.200  10.100 25.200  10.100 
      20.600  10.300 20.600  10.300 18.500  5.300 18.500  5.300 20.600  5.500 
      20.600  5.500 25.200  4.100 25.200  4.100 20.600  4.300 20.600  4.300 
      17.500  13.300 17.500  13.300 10.500  10.300 10.500  ;
      RECT 9.800 23.500  11.800 25.500  ;
      RECT 9.800 21.500  11.800 23.500  ;
      RECT 9.800 19.500  11.800 21.500  ;
      RECT 9.800 2.700  11.800 4.700  ;
      POLYGON 10.000 12.500  10.000 14.500  12.000 14.500  12.000 12.500  
      10.000 12.500  ;
      RECT 10.000 12.500  12.000 14.500  ;
      RECT 12.800 2.700  14.800 4.700  ;
      RECT 12.800 19.500  14.800 21.500  ;
      RECT 12.800 21.500  14.800 23.500  ;
      RECT 12.800 23.500  14.800 25.500  ;
      POLYGON 13.300 8.500  13.300 3.200  14.300 3.200  14.300 7.500  17.300 
      7.500  17.300 12.700  18.000 12.700  18.000 14.700  17.300 14.700  
      17.300 20.600  17.500 20.600  17.500 25.200  16.100 25.200  16.100 
      20.600  16.300 20.600  16.300 14.700  16.000 14.700  16.000 12.700  
      16.300 12.700  16.300 8.500  13.300 8.500  ;
      RECT 15.800 23.500  17.800 25.500  ;
      RECT 15.800 21.500  17.800 23.500  ;
      RECT 15.800 19.500  17.800 21.500  ;
    LAYER ML2 ;
      POLYGON 4.000 14.500  4.000 12.500  6.000 12.500  6.000 14.500  4.000 
      14.500  ;
      POLYGON 10.000 12.500  10.000 14.500  12.000 14.500  12.000 12.500  
      10.000 12.500  ;
      POLYGON 7.000 9.700  7.000 11.700  9.000 11.700  9.000 9.700  7.000 
      9.700  ;
      POLYGON 16.000 12.700  16.000 14.700  18.000 14.700  18.000 12.700  
      16.000 12.700  ;
      POLYGON 1.000 15.500  1.000 17.500  3.000 17.500  3.000 15.500  1.000 
      15.500  ;
    LAYER POL ;
      POLYGON 1.000 17.500  1.000 15.500  2.000 15.500  2.000 6.500  2.800 
      6.500  2.800 1.700  3.800 1.700  3.800 7.500  3.000 7.500  3.000 15.500  
      3.800 15.500  3.800 26.500  2.800 26.500  2.800 17.500  1.000 17.500  ;
      POLYGON 4.000 14.500  4.000 12.500  4.800 12.500  4.800 1.700  5.800 
      1.700  5.800 12.500  6.000 12.500  6.000 13.500  6.800 13.500  6.800 
      26.500  5.800 26.500  5.800 14.500  4.000 14.500  ;
      POLYGON 6.800 11.500  6.800 1.700  7.800 1.700  7.800 9.700  9.000 9.700 
       9.000 11.700  8.800 11.700  8.800 16.500  9.800 16.500  9.800 26.500  
      8.800 26.500  8.800 17.500  7.800 17.500  7.800 11.700  7.000 11.700  
      7.000 11.500  6.800 11.500  ;
      POLYGON 8.800 8.700  8.800 1.700  9.800 1.700  9.800 7.700  11.300 7.700 
       11.300 12.500  12.000 12.500  12.000 13.000  12.800 13.000  12.800 
      26.500  11.800 26.500  11.800 14.500  10.000 14.500  10.000 12.500  
      10.300 12.500  10.300 8.700  8.800 8.700  ;
      POLYGON 11.800 6.700  11.800 1.700  12.800 1.700  12.800 5.700  15.800 
      5.700  15.800 26.500  14.800 26.500  14.800 11.500  13.300 11.500  
      13.300 9.500  14.800 9.500  14.800 6.700  11.800 6.700  ;
    LAYER VIA1 ;
      POLYGON 10.500 13.000  10.500 14.000  11.500 14.000  11.500 13.000  
      10.500 13.000  ;
      POLYGON 7.500 10.200  7.500 11.200  8.500 11.200  8.500 10.200  7.500 
      10.200  ;
      POLYGON 4.500 13.000  4.500 14.000  5.500 14.000  5.500 13.000  4.500 
      13.000  ;
      POLYGON 16.500 13.200  16.500 14.200  17.500 14.200  17.500 13.200  
      16.500 13.200  ;
      POLYGON 1.500 16.000  1.500 17.000  2.500 17.000  2.500 16.000  1.500 
      16.000  ;
  END
END an41LEF


END LIBRARY
