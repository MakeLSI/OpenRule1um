VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO an21
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 12.500 BY 30.000 ;
  SYMMETRY X Y ;
  SITE unit ;
 
  PIN A
    USE SIGNAL ;
    PORT
      LAYER ML2 ;
        POLYGON 1.000 9.700  1.000 11.700  3.000 11.700  3.000 9.700  1.000 
        9.700  ;
    END
    PORT
      LAYER ML1 ;
        POLYGON 1.000 9.700  1.000 11.700  3.000 11.700  3.000 9.700  1.000 
        9.700  ;
    END
  END A
  PIN B
    USE SIGNAL ;
    PORT
      LAYER ML2 ;
        POLYGON 4.000 12.500  4.000 14.500  6.000 14.500  6.000 12.500  4.000 
        12.500  ;
    END
    PORT
      LAYER ML1 ;
        POLYGON 4.000 12.500  4.000 14.500  6.000 14.500  6.000 12.500  4.000 
        12.500  ;
    END
  END B
  PIN VDD
    USE POWER ;
    PORT
      LAYER ML1 ;
        RECT -0.500 28.500  13.000 30.500  ;
    END
  END VDD
  PIN VSS
    USE GROUND ;
    PORT
      LAYER ML1 ;
        RECT -0.500 -0.500  13.000 1.500  ;
    END
  END VSS
  PIN Y
    USE SIGNAL ;
    PORT
      LAYER ML2 ;
        POLYGON 10.000 12.500  10.000 14.500  12.000 14.500  12.000 12.500  
        10.000 12.500  ;
    END
    PORT
      LAYER ML1 ;
        POLYGON 10.000 12.500  10.000 14.500  12.000 14.500  12.000 12.500  
        10.000 12.500  ;
    END
    PORT
      LAYER ML1 ;
        WIDTH 1.000  ;
        PATH 10.800 20.500 10.800 6.500 9.800 6.500 9.800 3.800  ;
    END
  END Y
  OBS
    LAYER ML1 ;
      WIDTH 1.400  ;
      PATH 7.800 21.300 7.800 28.500  ;
      WIDTH 1.400  ;
      PATH 10.800 21.300 10.800 24.500  ;
      WIDTH 1.000  ;
      PATH 6.800 1.000 6.800 3.800  ;
      WIDTH 1.000  ;
      PATH 4.800 20.500 4.800 18.000 7.800 18.000 7.800 10.500 4.500 10.500 
      4.500 8.200 1.800 8.200 1.800 3.800  ;
      WIDTH 1.400  ;
      PATH 1.800 21.300 1.800 28.500  ;
      WIDTH 1.400  ;
      PATH 4.800 21.300 4.800 24.500  ;
    VIA 1.800 22.500  dcont ;
    VIA 1.800 20.500  dcont ;
    VIA 1.800 3.800  dcont ;
    VIA 1.800 24.500  dcont ;
    VIA 4.800 22.500  dcont ;
    VIA 4.800 20.500  dcont ;
    VIA 4.800 24.500  dcont ;
    VIA 6.800 3.800  dcont ;
    VIA 7.800 24.500  dcont ;
    VIA 7.800 22.500  dcont ;
    VIA 7.800 20.500  dcont ;
    VIA 9.800 3.800  dcont ;
    VIA 10.800 20.500  dcont ;
    VIA 10.800 22.500  dcont ;
    VIA 10.800 24.500  dcont ;
    VIA 5.000 13.500  pcont ;
    VIA 5.500 29.500  nsubcont ;
    VIA 8.300 10.500  pcont ;
    VIA 2.000 10.700  pcont ;
    VIA 5.000 0.500  psubcont ;
  END
END an21

MACRO dcont
  CLASS CORE ;
  OBS
    LAYER ML1 ;
      RECT -1.000 -1.000  1.000 1.000  ;
  END
END dcont

MACRO pcont
  CLASS CORE ;
  OBS
    LAYER ML1 ;
      RECT -1.000 -1.000  1.000 1.000  ;
  END
END pcont

MACRO nsubcont
  CLASS CORE ;
  OBS
    LAYER ML1 ;
      RECT -1.000 -1.000  1.000 1.000  ;
  END
END nsubcont

MACRO psubcont
  CLASS CORE ;
  OBS
    LAYER ML1 ;
      RECT -1.000 -1.000  1.000 1.000  ;
  END
END psubcont


END LIBRARY
