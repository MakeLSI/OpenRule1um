*******************************************************************************
* CDL netlist
*
* Library : OpenRule1um_StdCell
* Top Cell Name: rff1m2_r
* View Name: extracted
* Netlist created: 07.4.2020 15:10:02
*******************************************************************************

*.SCALE METER
*.GLOBAL vdd gnd

*******************************************************************************
* Library Name: OpenRule1um_StdCell
* Cell Name:    rff1m2_r
* View Name:    extracted
*******************************************************************************

.SUBCKT rff1m2_r

MM100 n15 n11 n1 n1 nch w=2e-06 l=1e-06 as=2e-12 ps=6e-06 ad=1e-12 pd=4e-06 $X=1.93e-05 $Y=2.8e-06
MM94 n1 n13 n12 n1 nch w=2e-06 l=1e-06 as=4e-12 ps=6e-06 ad=4e-12 pd=6e-06 $X=-3.7e-06 $Y=2.8e-06
MM95 n9 n12 n1 n1 nch w=2e-06 l=1e-06 as=4e-12 ps=6e-06 ad=4e-12 pd=6e-06 $X=2.8e-06 $Y=2.8e-06
MM109 n5 n4 n1 n1 nch w=2e-06 l=1e-06 as=4e-12 ps=6e-06 ad=4e-12 pd=6e-06 $X=4.93e-05 $Y=2.8e-06
MM113 n2 n9 n7 n2 pch w=6e-06 l=1e-06 as=6e-12 ps=1e-05 ad=6e-12 pd=1e-05 $X=5.8e-06 $Y=2.08e-05
MM110 n1 n5 n8 n1 nch w=2e-06 l=1e-06 as=2e-12 ps=6e-06 ad=2e-12 pd=6e-06 $X=5.23e-05 $Y=2.8e-06
MM122 n0 n9 n22 n2 pch w=6e-06 l=1e-06 as=3e-12 ps=8e-06 ad=6e-12 pd=1e-05 $X=3.58e-05 $Y=2.08e-05
MM125 n23 n3 n4 n2 pch w=6e-06 l=1e-06 as=6e-12 ps=1e-05 ad=3e-12 pd=8e-06 $X=4.28e-05 $Y=2.08e-05
MM112 n9 n12 n2 n2 pch w=6e-06 l=1e-06 as=1.2e-11 ps=1e-05 ad=1.2e-11 pd=1e-05 $X=2.8e-06 $Y=2.08e-05
MM126 n5 n4 n2 n2 pch w=6e-06 l=1e-06 as=1.2e-11 ps=1e-05 ad=1.2e-11 pd=1e-05 $X=4.93e-05 $Y=2.08e-05
MM108 n4 n3 n1 n1 nch w=2e-06 l=1e-06 as=1.9e-12 ps=5.8e-06 ad=2e-12 pd=6e-06 $X=4.13e-05 $Y=2.8e-06
MM99 n6 n9 n15 n1 nch w=2e-06 l=1e-06 as=1e-12 ps=4e-06 ad=2e-12 pd=6e-06 $X=1.73e-05 $Y=2.8e-06
MM97 n1 n10 n14 n1 nch w=2e-06 l=1e-06 as=2e-12 ps=4e-06 ad=4e-12 pd=6e-06 $X=1.23e-05 $Y=2.8e-06
MM115 n18 n9 n6 n2 pch w=6e-06 l=1e-06 as=6e-12 ps=1e-05 ad=3e-12 pd=8e-06 $X=1.43e-05 $Y=2.08e-05
MM103 n1 n11 n16 n1 nch w=2e-06 l=1e-06 as=1e-12 ps=4e-06 ad=2e-12 pd=6e-06 $X=2.83e-05 $Y=2.8e-06
MM111 n2 n13 n12 n2 pch w=6e-06 l=1e-06 as=1.2e-11 ps=1e-05 ad=1.2e-11 pd=1e-05 $X=-3.7e-06 $Y=1.95e-05
MM118 n2 n6 n20 n2 pch w=6e-06 l=1e-06 as=3e-12 ps=8e-06 ad=6e-12 pd=1e-05 $X=2.23e-05 $Y=2.08e-05
MM102 n11 n3 n1 n1 nch w=2e-06 l=1e-06 as=2e-12 ps=6e-06 ad=2e-12 pd=6e-06 $X=2.53e-05 $Y=2.8e-06
MM106 n17 n4 n1 n1 nch w=2e-06 l=1e-06 as=2e-12 ps=6e-06 ad=1e-12 pd=4e-06 $X=3.53e-05 $Y=2.8e-06
MM104 n16 n9 n0 n1 nch w=2e-06 l=1e-06 as=2e-12 ps=6e-06 ad=1e-12 pd=4e-06 $X=3.03e-05 $Y=2.8e-06
MM124 n2 n0 n23 n2 pch w=6e-06 l=1e-06 as=3e-12 ps=8e-06 ad=6e-12 pd=1e-05 $X=4.08e-05 $Y=2.08e-05
MM107 n1 n0 n4 n1 nch w=2e-06 l=1e-06 as=2e-12 ps=6e-06 ad=2e-12 pd=6e-06 $X=3.83e-05 $Y=2.8e-06
MM105 n0 n7 n17 n1 nch w=2e-06 l=1e-06 as=1e-12 ps=4e-06 ad=2e-12 pd=6e-06 $X=3.33e-05 $Y=2.8e-06
MM98 n14 n7 n6 n1 nch w=2e-06 l=1e-06 as=2e-12 ps=6e-06 ad=1e-12 pd=4e-06 $X=1.43e-05 $Y=2.8e-06
MM119 n20 n3 n11 n2 pch w=6e-06 l=1e-06 as=6e-12 ps=1e-05 ad=3e-12 pd=8e-06 $X=2.43e-05 $Y=2.08e-05
MM117 n19 n11 n2 n2 pch w=6e-06 l=1e-06 as=6e-12 ps=1e-05 ad=3e-12 pd=8e-06 $X=1.93e-05 $Y=2.08e-05
MM101 n1 n6 n11 n1 nch w=2e-06 l=1e-06 as=2e-12 ps=6e-06 ad=2e-12 pd=6e-06 $X=2.23e-05 $Y=2.8e-06
MM96 n1 n9 n7 n1 nch w=2e-06 l=1e-06 as=2e-12 ps=6e-06 ad=2e-12 pd=6e-06 $X=5.8e-06 $Y=2.8e-06
MM127 n2 n5 n8 n2 pch w=6e-06 l=1e-06 as=6e-12 ps=1e-05 ad=6e-12 pd=1e-05 $X=5.23e-05 $Y=2.08e-05
MM121 n21 n7 n0 n2 pch w=6e-06 l=1e-06 as=6e-12 ps=1e-05 ad=3e-12 pd=8e-06 $X=3.28e-05 $Y=2.08e-05
MM116 n6 n7 n19 n2 pch w=6e-06 l=1e-06 as=3e-12 ps=8e-06 ad=6e-12 pd=1e-05 $X=1.73e-05 $Y=2.08e-05
MM120 n2 n11 n21 n2 pch w=6e-06 l=1e-06 as=6e-12 ps=8e-06 ad=1.2e-11 pd=1e-05 $X=3.08e-05 $Y=2.08e-05
MM123 n22 n4 n2 n2 pch w=6e-06 l=1e-06 as=6e-12 ps=1e-05 ad=3e-12 pd=8e-06 $X=3.78e-05 $Y=2.08e-05
MM114 n2 n10 n18 n2 pch w=6e-06 l=1e-06 as=6e-12 ps=8e-06 ad=1.2e-11 pd=1e-05 $X=1.23e-05 $Y=2.08e-05
.ENDS
