VERSION 5.3 ;

NAMESCASESENSITIVE ON ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS











MACRO buf4LEF
  CLASS BLOCK ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER ML1 ;
        POLYGON 1.000 14.500  1.000 16.500  3.000 16.500  3.000 14.500  1.000 
        14.500  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    PORT
      LAYER ML1 ;
        POLYGON -0.500 30.500  -0.500 28.500  4.100 28.500  4.100 20.600  
        5.500 20.600  5.500 28.500  10.100 28.500  10.100 20.600  11.500 
        20.600  11.500 28.500  16.100 28.500  16.100 20.600  17.500 20.600  
        17.500 28.500  19.000 28.500  19.000 30.500  -0.500 30.500  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    PORT
      LAYER ML1 ;
        POLYGON -0.500 1.500  -0.500 -0.500  19.000 -0.500  19.000 1.500  
        17.300 1.500  17.300 4.200  16.300 4.200  16.300 1.500  11.300 1.500  
        11.300 4.200  10.300 4.200  10.300 1.500  5.300 1.500  5.300 4.200  
        4.300 4.200  4.300 1.500  -0.500 1.500  ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    PORT
      LAYER ML1 ;
        POLYGON 7.100 25.200  7.100 20.600  7.300 20.600  7.300 3.300  8.300 
        3.300  8.300 7.000  13.300 7.000  13.300 3.300  14.300 3.300  14.300 
        15.000  15.000 15.000  15.000 17.000  14.300 17.000  14.300 20.600  
        14.500 20.600  14.500 25.200  13.100 25.200  13.100 20.600  13.300 
        20.600  13.300 17.000  13.000 17.000  13.000 15.000  13.300 15.000  
        13.300 9.000  8.300 9.000  8.300 20.600  8.500 20.600  8.500 25.200  
        7.100 25.200  ;
    END
  END Y
  OBS
    LAYER CNT ;
      POLYGON 13.300 22.000  13.300 23.000  14.300 23.000  14.300 22.000  
      13.300 22.000  ;
      POLYGON 13.300 24.000  13.300 25.000  14.300 25.000  14.300 24.000  
      13.300 24.000  ;
      POLYGON 13.300 3.200  13.300 4.200  14.300 4.200  14.300 3.200  13.300 
      3.200  ;
      POLYGON 16.300 20.000  16.300 21.000  17.300 21.000  17.300 20.000  
      16.300 20.000  ;
      POLYGON 16.300 22.000  16.300 23.000  17.300 23.000  17.300 22.000  
      16.300 22.000  ;
      POLYGON 16.300 24.000  16.300 25.000  17.300 25.000  17.300 24.000  
      16.300 24.000  ;
      POLYGON 16.300 3.200  16.300 4.200  17.300 4.200  17.300 3.200  16.300 
      3.200  ;
      POLYGON 4.800 11.000  4.800 12.000  5.800 12.000  5.800 11.000  4.800 
      11.000  ;
      POLYGON 4.500 29.000  4.500 30.000  5.500 30.000  5.500 29.000  4.500 
      29.000  ;
      POLYGON 1.500 15.000  1.500 16.000  2.500 16.000  2.500 15.000  1.500 
      15.000  ;
      POLYGON 4.500 0.000  4.500 1.000  5.500 1.000  5.500 0.000  4.500 0.000  ;
      
      POLYGON 13.300 20.000  13.300 21.000  14.300 21.000  14.300 20.000  
      13.300 20.000  ;
      POLYGON 10.300 24.000  10.300 25.000  11.300 25.000  11.300 24.000  
      10.300 24.000  ;
      POLYGON 10.300 22.000  10.300 23.000  11.300 23.000  11.300 22.000  
      10.300 22.000  ;
      POLYGON 10.300 20.000  10.300 21.000  11.300 21.000  11.300 20.000  
      10.300 20.000  ;
      POLYGON 10.300 3.200  10.300 4.200  11.300 4.200  11.300 3.200  10.300 
      3.200  ;
      POLYGON 7.300 3.200  7.300 4.200  8.300 4.200  8.300 3.200  7.300 3.200  ;
      
      POLYGON 7.300 20.000  7.300 21.000  8.300 21.000  8.300 20.000  7.300 
      20.000  ;
      POLYGON 7.300 22.000  7.300 23.000  8.300 23.000  8.300 22.000  7.300 
      22.000  ;
      POLYGON 7.300 24.000  7.300 25.000  8.300 25.000  8.300 24.000  7.300 
      24.000  ;
      POLYGON 4.300 22.000  4.300 23.000  5.300 23.000  5.300 22.000  4.300 
      22.000  ;
      POLYGON 4.300 20.000  4.300 21.000  5.300 21.000  5.300 20.000  4.300 
      20.000  ;
      POLYGON 4.300 24.000  4.300 25.000  5.300 25.000  5.300 24.000  4.300 
      24.000  ;
      POLYGON 4.300 3.200  4.300 4.200  5.300 4.200  5.300 3.200  4.300 3.200  ;
      
      POLYGON 1.300 22.000  1.300 23.000  2.300 23.000  2.300 22.000  1.300 
      22.000  ;
      POLYGON 1.300 20.000  1.300 21.000  2.300 21.000  2.300 20.000  1.300 
      20.000  ;
      POLYGON 1.300 3.200  1.300 4.200  2.300 4.200  2.300 3.200  1.300 3.200  ;
      
      POLYGON 1.300 24.000  1.300 25.000  2.300 25.000  2.300 24.000  1.300 
      24.000  ;
    LAYER FRAME ;
      POLYGON -0.500 1.500  -0.500 -0.500  19.000 -0.500  19.000 1.500  -0.500 
      1.500  ;
      POLYGON 0.000 0.000  18.500 0.000  18.500 30.000  0.000 30.000  0.000 
      0.000  ;
      RECT -0.500 28.500  19.000 30.500  ;
    LAYER ML1 ;
      WIDTH 1.400  ;
      PATH 10.800 21.300 10.800 24.500  ;
      POLYGON 1.000 14.500  1.000 16.500  3.000 16.500  3.000 14.500  1.000 
      14.500  ;
      RECT 4.000 -0.500  6.000 1.500  ;
      RECT 1.000 14.500  3.000 16.500  ;
      RECT 4.000 28.500  6.000 30.500  ;
      RECT 15.800 2.700  17.800 4.700  ;
      RECT 15.800 23.500  17.800 25.500  ;
      RECT 15.800 21.500  17.800 23.500  ;
      RECT 15.800 19.500  17.800 21.500  ;
      RECT 12.800 2.700  14.800 4.700  ;
      RECT 12.800 23.500  14.800 25.500  ;
      RECT 12.800 21.500  14.800 23.500  ;
      RECT 12.800 19.500  14.800 21.500  ;
      RECT 9.800 23.500  11.800 25.500  ;
      RECT 9.800 21.500  11.800 23.500  ;
      RECT 9.800 19.500  11.800 21.500  ;
      RECT 9.800 2.700  11.800 4.700  ;
      RECT 6.800 2.700  8.800 4.700  ;
      RECT 6.800 19.500  8.800 21.500  ;
      RECT 6.800 21.500  8.800 23.500  ;
      RECT 6.800 23.500  8.800 25.500  ;
      RECT 3.800 21.500  5.800 23.500  ;
      RECT 3.800 19.500  5.800 21.500  ;
      RECT 3.800 23.500  5.800 25.500  ;
      RECT 3.800 2.700  5.800 4.700  ;
      RECT 0.800 21.500  2.800 23.500  ;
      RECT 0.800 19.500  2.800 21.500  ;
      RECT 0.800 2.700  2.800 4.700  ;
      RECT 0.800 23.500  2.800 25.500  ;
      POLYGON -0.500 30.500  -0.500 28.500  4.100 28.500  4.100 20.600  5.500 
      20.600  5.500 28.500  10.100 28.500  10.100 20.600  11.500 20.600  
      11.500 28.500  16.100 28.500  16.100 20.600  17.500 20.600  17.500 
      28.500  19.000 28.500  19.000 30.500  -0.500 30.500  ;
      POLYGON 1.300 8.000  1.300 3.200  2.300 3.200  2.300 7.000  5.000 7.000  
      5.000 10.500  6.300 10.500  6.300 12.500  5.000 12.500  5.000 18.500  
      2.300 18.500  2.300 20.600  2.500 20.600  2.500 25.200  1.100 25.200  
      1.100 20.600  1.300 20.600  1.300 17.500  4.000 17.500  4.000 8.000  
      1.300 8.000  ;
      POLYGON 7.100 25.200  7.100 20.600  7.300 20.600  7.300 3.300  8.300 
      3.300  8.300 7.000  13.300 7.000  13.300 3.300  14.300 3.300  14.300 
      15.000  15.000 15.000  15.000 17.000  14.300 17.000  14.300 20.600  
      14.500 20.600  14.500 25.200  13.100 25.200  13.100 20.600  13.300 
      20.600  13.300 17.000  13.000 17.000  13.000 15.000  13.300 15.000  
      13.300 9.000  8.300 9.000  8.300 20.600  8.500 20.600  8.500 25.200  
      7.100 25.200  ;
      POLYGON -0.500 1.500  -0.500 -0.500  19.000 -0.500  19.000 1.500  17.300 
      1.500  17.300 4.200  16.300 4.200  16.300 1.500  11.300 1.500  11.300 
      4.200  10.300 4.200  10.300 1.500  5.300 1.500  5.300 4.200  4.300 4.200 
       4.300 1.500  -0.500 1.500  ;
    LAYER ML2 ;
      POLYGON 13.000 15.000  13.000 17.000  15.000 17.000  15.000 15.000  
      13.000 15.000  ;
      POLYGON 1.000 14.500  1.000 16.500  3.000 16.500  3.000 14.500  1.000 
      14.500  ;
    LAYER POL ;
      POLYGON 4.300 12.500  4.300 10.500  5.800 10.500  5.800 1.700  6.800 
      1.700  6.800 10.500  8.800 10.500  8.800 1.700  9.800 1.700  9.800 
      10.500  11.800 10.500  11.800 1.700  12.800 1.700  12.800 10.500  14.800 
      10.500  14.800 1.700  15.800 1.700  15.800 26.500  14.800 26.500  14.800 
      12.500  12.800 12.500  12.800 26.500  11.800 26.500  11.800 12.500  
      9.800 12.500  9.800 26.500  8.800 26.500  8.800 12.500  6.800 12.500  
      6.800 26.500  5.800 26.500  5.800 12.500  4.300 12.500  ;
      POLYGON 1.000 16.500  1.000 14.500  1.500 14.500  1.500 8.500  2.800 
      8.500  2.800 1.700  3.800 1.700  3.800 9.500  2.500 9.500  2.500 14.500  
      3.000 14.500  3.000 15.500  3.800 15.500  3.800 26.500  2.800 26.500  
      2.800 16.500  1.000 16.500  ;
    LAYER VIA1 ;
      POLYGON 13.500 15.500  13.500 16.500  14.500 16.500  14.500 15.500  
      13.500 15.500  ;
      POLYGON 1.500 15.000  1.500 16.000  2.500 16.000  2.500 15.000  1.500 
      15.000  ;
  END
END buf4LEF


END LIBRARY
