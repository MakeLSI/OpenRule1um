*******************************************************************************
* CDL netlist
*
* Library : OpenRule1um_StdCell
* Top Cell Name: sff1_r
* View Name: schematic
* Netlist created: 07.4.2020 15:15:01
*******************************************************************************

*.SCALE METER
*.GLOBAL VDD VSS

*******************************************************************************
* Library Name: OpenRule1um_StdCell
* Cell Name:    sff1_r
* View Name:    schematic
*******************************************************************************

.SUBCKT sff1_r CK S Q D 
*.PININFO CK:I S:I Q:O D:I QB:O

M24 n8 n5 n9 VDD pch w=6u l=1u m=1
M20 n9 n5 n10 VSS nch w=2u l=1u m=1
M29 n23 n9 VSS VSS nch w=2u l=1u m=1
M2 n16 n13 n11 VDD pch w=6u l=1u m=1
M26 n9 n13 n21 VSS nch w=2u l=1u m=1
M27 n10 n7 VSS VSS nch w=2u l=1u m=1
M22 VDD n7 n22 VDD pch w=6u l=1u m=1
M0 VDD n13 n5 VDD pch w=6u l=1u m=1
M14 VDD S n3 VDD pch w=6u l=1u m=1
M12 VDD n11 n3 VDD pch w=6u l=1u m=1
M4 n11 n5 n15 VSS nch w=2u l=1u m=1
M6 n13 n25 VSS VSS nch w=2u l=1u m=1
M17 VDD S n7 VDD pch w=6u l=1u m=1
M28 n7 S n23 VSS nch w=2u l=1u m=1
M23 n21 n3 VSS VSS nch w=2u l=1u m=1
M19 VDD n9 n7 VDD pch w=6u l=1u m=1
M11 n11 n13 n20 VSS nch w=2u l=1u m=1
M16 n12 n11 VSS VSS nch w=2u l=1u m=1
M9 n20 n3 VSS VSS nch w=2u l=1u m=1
M15 n3 S n12 VSS nch w=2u l=1u m=1
M34 n25 CK VSS VSS nch w=2u l=1u m=1
M30 VDD n7 QB VDD pch w=6u l=1u m=1
M25 VDD n3 n8 VDD pch w=6u l=1u m=1
M5 n15 D VSS VSS nch w=2u l=1u m=1
M32_40 Q QB VSS VSS nch w=2u l=1u m=1
M21 n22 n13 n9 VDD pch w=6u l=1u m=1
M3 VDD D n16 VDD pch w=6u l=1u m=1
M8 VDD n3 n14 VDD pch w=6u l=1u m=1
M7 VDD n25 n13 VDD pch w=6u l=1u m=1
M32 VDD CK n25 VDD pch w=6u l=1u m=1
M31 VDD QB Q VDD pch w=6u l=1u m=1
M1 n5 n13 VSS VSS nch w=2u l=1u m=1
M10 n14 n5 n11 VDD pch w=6u l=1u m=1
M33 QB n7 VSS VSS nch w=2u l=1u m=1
.ENDS

