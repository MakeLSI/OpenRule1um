VERSION 5.3 ;

NAMESCASESENSITIVE ON ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS











MACRO nr222LEF
  CLASS BLOCK ;
  PIN A0
    DIRECTION INPUT ;
    PORT
      LAYER POL ;
        POLYGON 1.000 16.500  1.000 14.500  2.000 14.500  2.000 6.000  2.800 
        6.000  2.800 1.700  3.800 1.700  3.800 7.000  3.000 7.000  3.000 
        15.000  3.800 15.000  3.800 26.500  2.800 26.500  2.800 16.500  1.000 
        16.500  ;
    END
    PORT
      LAYER ML1 ;
        POLYGON 1.000 14.500  1.000 16.500  3.000 16.500  3.000 14.500  1.000 
        14.500  ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER POL ;
        POLYGON 4.000 10.500  4.000 8.500  4.800 8.500  4.800 1.700  5.800 
        1.700  5.800 8.500  6.000 8.500  6.000 15.000  6.800 15.000  6.800 
        26.500  5.800 26.500  5.800 16.000  5.000 16.000  5.000 10.500  4.000 
        10.500  ;
    END
    PORT
      LAYER ML1 ;
        POLYGON 4.000 8.500  4.000 10.500  6.000 10.500  6.000 8.500  4.000 
        8.500  ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    PORT
      LAYER POL ;
        POLYGON 9.800 8.500  9.800 1.700  10.800 1.700  10.800 7.500  12.800 
        7.500  12.800 26.500  11.800 26.500  11.800 16.500  10.000 16.500  
        10.000 14.500  11.800 14.500  11.800 8.500  9.800 8.500  ;
    END
    PORT
      LAYER ML1 ;
        POLYGON 10.000 14.500  10.000 16.500  12.000 16.500  12.000 14.500  
        10.000 14.500  ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER POL ;
        POLYGON 7.000 13.500  7.000 11.500  7.800 11.500  7.800 1.700  8.800 
        1.700  8.800 11.500  9.000 11.500  9.000 17.500  9.800 17.500  9.800 
        26.500  8.800 26.500  8.800 18.500  8.000 18.500  8.000 13.500  7.000 
        13.500  ;
    END
    PORT
      LAYER ML1 ;
        POLYGON 7.000 11.500  7.000 13.500  9.000 13.500  9.000 11.500  7.000 
        11.500  ;
    END
  END B1
  PIN VDD
    DIRECTION INOUT ;
    PORT
      LAYER ML1 ;
        POLYGON -0.500 30.500  -0.500 28.500  4.100 28.500  4.100 20.600  
        5.500 20.600  5.500 28.500  16.000 28.500  16.000 30.500  -0.500 
        30.500  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    PORT
      LAYER ML1 ;
        POLYGON -0.500 1.500  -0.500 -0.500  16.000 -0.500  16.000 1.500  
        12.300 1.500  12.300 4.200  11.300 4.200  11.300 1.500  2.300 1.500  
        2.300 4.200  1.300 4.200  1.300 1.500  -0.500 1.500  ;
    END
  END VSS
  PIN YB
    DIRECTION OUTPUT ;
    PORT
      LAYER ML1 ;
        POLYGON 6.300 7.000  6.300 3.200  7.300 3.200  7.300 6.000  14.000 
        6.000  14.000 8.000  14.500 8.000  14.500 10.000  14.000 10.000  
        14.000 18.500  11.300 18.500  11.300 20.600  11.500 20.600  11.500 
        25.200  10.100 25.200  10.100 20.600  10.300 20.600  10.300 17.500  
        13.000 17.500  13.000 10.000  12.500 10.000  12.500 8.000  13.000 
        8.000  13.000 7.000  6.300 7.000  ;
    END
  END YB
  OBS
    LAYER CNT ;
      POLYGON 10.300 24.000  10.300 25.000  11.300 25.000  11.300 24.000  
      10.300 24.000  ;
      POLYGON 11.300 3.200  11.300 4.200  12.300 4.200  12.300 3.200  11.300 
      3.200  ;
      POLYGON 13.300 20.000  13.300 21.000  14.300 21.000  14.300 20.000  
      13.300 20.000  ;
      POLYGON 13.300 22.000  13.300 23.000  14.300 23.000  14.300 22.000  
      13.300 22.000  ;
      POLYGON 13.300 24.000  13.300 25.000  14.300 25.000  14.300 24.000  
      13.300 24.000  ;
      POLYGON 10.500 15.000  10.500 16.000  11.500 16.000  11.500 15.000  
      10.500 15.000  ;
      POLYGON 7.500 12.000  7.500 13.000  8.500 13.000  8.500 12.000  7.500 
      12.000  ;
      POLYGON 9.700 29.000  9.700 30.000  10.700 30.000  10.700 29.000  9.700 
      29.000  ;
      POLYGON 4.500 9.000  4.500 10.000  5.500 10.000  5.500 9.000  4.500 
      9.000  ;
      POLYGON 1.500 15.000  1.500 16.000  2.500 16.000  2.500 15.000  1.500 
      15.000  ;
      POLYGON 9.700 0.000  9.700 1.000  10.700 1.000  10.700 0.000  9.700 
      0.000  ;
      POLYGON 10.300 22.000  10.300 23.000  11.300 23.000  11.300 22.000  
      10.300 22.000  ;
      POLYGON 10.300 20.000  10.300 21.000  11.300 21.000  11.300 20.000  
      10.300 20.000  ;
      POLYGON 7.300 20.000  7.300 21.000  8.300 21.000  8.300 20.000  7.300 
      20.000  ;
      POLYGON 7.300 22.000  7.300 23.000  8.300 23.000  8.300 22.000  7.300 
      22.000  ;
      POLYGON 7.300 24.000  7.300 25.000  8.300 25.000  8.300 24.000  7.300 
      24.000  ;
      POLYGON 6.300 3.200  6.300 4.200  7.300 4.200  7.300 3.200  6.300 3.200  ;
      
      POLYGON 4.300 24.000  4.300 25.000  5.300 25.000  5.300 24.000  4.300 
      24.000  ;
      POLYGON 4.300 20.000  4.300 21.000  5.300 21.000  5.300 20.000  4.300 
      20.000  ;
      POLYGON 4.300 22.000  4.300 23.000  5.300 23.000  5.300 22.000  4.300 
      22.000  ;
      POLYGON 1.300 24.000  1.300 25.000  2.300 25.000  2.300 24.000  1.300 
      24.000  ;
      POLYGON 1.300 3.200  1.300 4.200  2.300 4.200  2.300 3.200  1.300 3.200  ;
      
      POLYGON 1.300 20.000  1.300 21.000  2.300 21.000  2.300 20.000  1.300 
      20.000  ;
      POLYGON 1.300 22.000  1.300 23.000  2.300 23.000  2.300 22.000  1.300 
      22.000  ;
    LAYER FRAME ;
      RECT -0.500 28.500  16.000 30.500  ;
      RECT -0.500 -0.500  16.000 1.500  ;
      POLYGON 0.000 0.000  15.500 0.000  15.500 30.000  0.000 30.000  0.000 
      0.000  ;
    LAYER ML1 ;
      POLYGON 1.000 14.500  1.000 16.500  3.000 16.500  3.000 14.500  1.000 
      14.500  ;
      WIDTH 1.400  ;
      PATH 1.800 21.300 1.800 24.500  ;
      POLYGON 4.000 8.500  4.000 10.500  6.000 10.500  6.000 8.500  4.000 
      8.500  ;
      RECT 9.200 -0.500  11.200 1.500  ;
      POLYGON 7.000 11.500  7.000 13.500  9.000 13.500  9.000 11.500  7.000 
      11.500  ;
      POLYGON 10.000 14.500  10.000 16.500  12.000 16.500  12.000 14.500  
      10.000 14.500  ;
      RECT 1.000 14.500  3.000 16.500  ;
      RECT 4.000 8.500  6.000 10.500  ;
      RECT 9.200 28.500  11.200 30.500  ;
      RECT 7.000 11.500  9.000 13.500  ;
      RECT 10.000 14.500  12.000 16.500  ;
      RECT 12.800 23.500  14.800 25.500  ;
      RECT 12.800 21.500  14.800 23.500  ;
      RECT 12.800 19.500  14.800 21.500  ;
      RECT 10.800 2.700  12.800 4.700  ;
      RECT 9.800 23.500  11.800 25.500  ;
      RECT 9.800 21.500  11.800 23.500  ;
      RECT 9.800 19.500  11.800 21.500  ;
      RECT 6.800 19.500  8.800 21.500  ;
      RECT 6.800 21.500  8.800 23.500  ;
      RECT 6.800 23.500  8.800 25.500  ;
      RECT 5.800 2.700  7.800 4.700  ;
      RECT 3.800 23.500  5.800 25.500  ;
      RECT 3.800 19.500  5.800 21.500  ;
      RECT 3.800 21.500  5.800 23.500  ;
      RECT 0.800 23.500  2.800 25.500  ;
      RECT 0.800 2.700  2.800 4.700  ;
      RECT 0.800 19.500  2.800 21.500  ;
      RECT 0.800 21.500  2.800 23.500  ;
      POLYGON -0.500 30.500  -0.500 28.500  4.100 28.500  4.100 20.600  5.500 
      20.600  5.500 28.500  16.000 28.500  16.000 30.500  -0.500 30.500  ;
      POLYGON -0.500 1.500  -0.500 -0.500  16.000 -0.500  16.000 1.500  12.300 
      1.500  12.300 4.200  11.300 4.200  11.300 1.500  2.300 1.500  2.300 
      4.200  1.300 4.200  1.300 1.500  -0.500 1.500  ;
      POLYGON 6.300 7.000  6.300 3.200  7.300 3.200  7.300 6.000  14.000 6.000 
       14.000 8.000  14.500 8.000  14.500 10.000  14.000 10.000  14.000 18.500 
       11.300 18.500  11.300 20.600  11.500 20.600  11.500 25.200  10.100 
      25.200  10.100 20.600  10.300 20.600  10.300 17.500  13.000 17.500  
      13.000 10.000  12.500 10.000  12.500 8.000  13.000 8.000  13.000 7.000  
      6.300 7.000  ;
      POLYGON 1.300 25.000  1.300 17.500  8.300 17.500  8.300 26.500  13.300 
      26.500  13.300 20.000  14.300 20.000  14.300 27.500  7.300 27.500  7.300 
      18.500  2.300 18.500  2.300 25.000  1.300 25.000  ;
    LAYER ML2 ;
      POLYGON 12.500 10.000  12.500 8.000  14.500 8.000  14.500 10.000  12.500 
      10.000  ;
      POLYGON 10.000 14.500  10.000 16.500  12.000 16.500  12.000 14.500  
      10.000 14.500  ;
      POLYGON 7.000 11.500  7.000 13.500  9.000 13.500  9.000 11.500  7.000 
      11.500  ;
      POLYGON 4.000 8.500  4.000 10.500  6.000 10.500  6.000 8.500  4.000 
      8.500  ;
      POLYGON 1.000 14.500  1.000 16.500  3.000 16.500  3.000 14.500  1.000 
      14.500  ;
    LAYER POL ;
      POLYGON 9.800 8.500  9.800 1.700  10.800 1.700  10.800 7.500  12.800 
      7.500  12.800 26.500  11.800 26.500  11.800 16.500  10.000 16.500  
      10.000 14.500  11.800 14.500  11.800 8.500  9.800 8.500  ;
      POLYGON 7.000 13.500  7.000 11.500  7.800 11.500  7.800 1.700  8.800 
      1.700  8.800 11.500  9.000 11.500  9.000 17.500  9.800 17.500  9.800 
      26.500  8.800 26.500  8.800 18.500  8.000 18.500  8.000 13.500  7.000 
      13.500  ;
      POLYGON 4.000 10.500  4.000 8.500  4.800 8.500  4.800 1.700  5.800 1.700 
       5.800 8.500  6.000 8.500  6.000 15.000  6.800 15.000  6.800 26.500  
      5.800 26.500  5.800 16.000  5.000 16.000  5.000 10.500  4.000 10.500  ;
      POLYGON 1.000 16.500  1.000 14.500  2.000 14.500  2.000 6.000  2.800 
      6.000  2.800 1.700  3.800 1.700  3.800 7.000  3.000 7.000  3.000 15.000  
      3.800 15.000  3.800 26.500  2.800 26.500  2.800 16.500  1.000 16.500  ;
    LAYER VIA1 ;
      POLYGON 10.500 15.000  10.500 16.000  11.500 16.000  11.500 15.000  
      10.500 15.000  ;
      POLYGON 7.500 12.000  7.500 13.000  8.500 13.000  8.500 12.000  7.500 
      12.000  ;
      POLYGON 4.500 9.000  4.500 10.000  5.500 10.000  5.500 9.000  4.500 
      9.000  ;
      POLYGON 13.000 8.500  13.000 9.500  14.000 9.500  14.000 8.500  13.000 
      8.500  ;
      POLYGON 1.500 15.000  1.500 16.000  2.500 16.000  2.500 15.000  1.500 
      15.000  ;
  END
END nr222LEF


END LIBRARY
