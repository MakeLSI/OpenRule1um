VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO inv8
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 27.500 BY 30.000 ;
  SYMMETRY X Y ;
  SITE unit ;
  
  PIN A
    USE SIGNAL ;
    PORT
      LAYER ML2 ;
        POLYGON 1.000 14.500  1.000 16.500  3.000 16.500  3.000 14.500  1.000 
        14.500  ;
    END
    PORT
      LAYER ML1 ;
        POLYGON 1.000 14.500  1.000 16.500  3.000 16.500  3.000 14.500  1.000 
        14.500  ;
    END
  END A
  PIN VDD
    USE POWER ;
    PORT
      LAYER ML1 ;
        RECT -0.500 28.500  28.000 30.500  ;
    END
  END VDD
  PIN VSS
    USE GROUND ;
    PORT
      LAYER ML1 ;
        RECT -0.500 -0.500  28.000 1.500  ;
    END
  END VSS
  PIN YB
    USE SIGNAL ;
    PORT
      LAYER ML1 ;
        WIDTH 1.000  ;
        PATH 4.800 11.000 22.800 11.000  ;
    END
    PORT
      LAYER ML1 ;
        WIDTH 1.000  ;
        PATH 4.800 20.500 4.800 3.800  ;
    END
    PORT
      LAYER ML1 ;
        WIDTH 1.000  ;
        PATH 10.800 20.500 10.800 3.800  ;
    END
    PORT
      LAYER ML1 ;
        WIDTH 1.000  ;
        PATH 16.800 20.500 16.800 3.800  ;
    END
    PORT
      LAYER ML1 ;
        POLYGON 22.000 10.500  22.000 12.500  24.000 12.500  24.000 10.500  
        22.000 10.500  ;
    END
    PORT
      LAYER ML2 ;
        POLYGON 22.000 10.500  22.000 12.500  24.000 12.500  24.000 10.500  
        22.000 10.500  ;
    END
    PORT
      LAYER ML1 ;
        WIDTH 1.000  ;
        PATH 22.800 20.500 22.800 3.800  ;
    END
  END YB
  OBS

    LAYER ML1 ;
      WIDTH 1.000  ;
      PATH 1.800 1.000 1.800 3.800  ;
      WIDTH 1.400  ;
      PATH 1.800 21.300 1.800 28.500  ;
      WIDTH 1.000  ;
      PATH 4.800 20.500 4.800 3.800  ;
      WIDTH 1.400  ;
      PATH 4.800 21.300 4.800 24.500  ;
      WIDTH 1.000  ;
      PATH 7.800 1.000 7.800 3.800  ;
      WIDTH 1.400  ;
      PATH 7.800 21.300 7.800 28.500  ;
      WIDTH 1.000  ;
      PATH 10.800 20.500 10.800 3.800  ;
      WIDTH 1.400  ;
      PATH 10.800 21.300 10.800 24.500  ;

      WIDTH 1.400  ;
      PATH 13.800 21.300 13.800 28.500  ;
      WIDTH 1.000  ;
      PATH 4.800 11.000 22.800 11.000  ;
      WIDTH 1.000  ;
      PATH 13.800 1.000 13.800 3.800  ;
      WIDTH 1.000  ;
      PATH 16.800 20.500 16.800 3.800  ;
      WIDTH 1.400  ;
      PATH 19.800 21.300 19.800 24.500  ;
      WIDTH 1.400  ;
      PATH 19.800 21.300 19.800 28.500  ;
      WIDTH 1.000  ;
      PATH 19.800 1.000 19.800 3.800  ;
      WIDTH 1.000  ;
      PATH 22.800 20.500 22.800 3.800  ;
      WIDTH 1.400  ;
      PATH 25.800 21.300 25.800 24.500  ;
      WIDTH 1.400  ;
      PATH 25.800 21.300 25.800 28.500  ;
      WIDTH 1.000  ;
      PATH 25.800 1.000 25.800 3.800  ;

    VIA 1.800 3.800  dcont ;
    VIA 1.800 22.500  dcont ;
    VIA 1.800 20.500  dcont ;
    VIA 1.800 24.500  dcont ;
    VIA 4.800 3.800  dcont ;
    VIA 4.800 22.500  dcont ;
    VIA 4.800 20.500  dcont ;
    VIA 4.800 24.500  dcont ;
    VIA 7.800 3.800  dcont ;
    VIA 7.800 20.500  dcont ;
    VIA 7.800 22.500  dcont ;
    VIA 7.800 24.500  dcont ;
    VIA 10.800 24.500  dcont ;
    VIA 10.800 20.500  dcont ;
    VIA 10.800 22.500  dcont ;
    VIA 10.800 3.800  dcont ;
    VIA 13.800 20.500  dcont ;
    VIA 13.800 22.500  dcont ;
    VIA 13.800 24.500  dcont ;
    VIA 13.800 3.800  dcont ;
    VIA 16.800 24.500  dcont ;
    VIA 16.800 20.500  dcont ;
    VIA 16.800 22.500  dcont ;
    VIA 16.800 3.800  dcont ;
    VIA 19.800 24.500  dcont ;
    VIA 19.800 20.500  dcont ;
    VIA 19.800 22.500  dcont ;
    VIA 19.800 3.800  dcont ;
    VIA 22.800 24.500  dcont ;
    VIA 22.800 22.500  dcont ;
    VIA 22.800 20.500  dcont ;
    VIA 22.800 3.800  dcont ;
    VIA 25.800 22.500  dcont ;
    VIA 25.800 20.500  dcont ;
    VIA 25.800 24.500  dcont ;
    VIA 25.800 3.800  dcont ;
    VIA 5.000 29.500  nsubcont ;
    VIA 18.300 0.500  psubcont ;
    VIA 2.000 15.500  pcont ;
    VIA 5.000 0.500  psubcont ;
    VIA 19.100 29.500  nsubcont ;
  END
END inv8

MACRO dcont
  CLASS CORE ;
  OBS
    LAYER ML1 ;
      RECT -1.000 -1.000  1.000 1.000  ;
  END
END dcont

MACRO nsubcont
  CLASS CORE ;
  OBS
    LAYER ML1 ;
      RECT -1.000 -1.000  1.000 1.000  ;
  END
END nsubcont

MACRO psubcont
  CLASS CORE ;
  OBS
    LAYER ML1 ;
      RECT -1.000 -1.000  1.000 1.000  ;
  END
END psubcont

MACRO pcont
  CLASS CORE ;
  OBS
    LAYER ML1 ;
      RECT -1.000 -1.000  1.000 1.000  ;
  END
END pcont


END LIBRARY
