VERSION 5.3 ;

NAMESCASESENSITIVE ON ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS











MACRO exorLEF
  CLASS BLOCK ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER POL ;
        POLYGON 5.800 8.000  5.800 1.700  6.800 1.700  6.800 7.000  7.000 
        7.000  7.000 13.700  8.000 13.700  8.000 15.700  7.000 15.700  7.000 
        18.000  5.800 18.000  5.800 27.800  4.800 27.800  4.800 17.000  6.000 
        17.000  6.000 8.000  5.800 8.000  ;
    END
    PORT
      LAYER ML1 ;
        RECT 6.000 13.700  8.000 15.700  ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER POL ;
        POLYGON 2.800 27.800  2.800 1.700  3.800 1.700  3.800 9.700  5.000 
        9.700  5.000 11.700  3.800 11.700  3.800 27.800  2.800 27.800  ;
    END
    PORT
      LAYER ML1 ;
        POLYGON 3.000 11.700  3.000 9.700  5.000 9.700  5.000 10.200  10.300 
        10.200  10.300 9.700  12.300 9.700  12.300 11.700  10.300 11.700  
        10.300 11.200  5.000 11.200  5.000 11.700  3.000 11.700  ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    PORT
      LAYER ML1 ;
        POLYGON -0.500 30.500  -0.500 28.500  6.100 28.500  6.100 21.900  
        7.500 21.900  7.500 28.500  12.600 28.500  12.600 21.900  14.000 
        21.900  14.000 28.500  21.500 28.500  21.500 30.500  -0.500 30.500  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    PORT
      LAYER ML1 ;
        POLYGON -0.500 1.500  -0.500 -0.500  21.500 -0.500  21.500 1.500  
        18.800 1.500  18.800 4.200  17.800 4.200  17.800 1.500  10.800 1.500  
        10.800 4.200  9.800 4.200  9.800 1.500  8.300 1.500  8.300 4.200  
        7.300 4.200  7.300 1.500  2.300 1.500  2.300 4.200  1.300 4.200  1.300 
        1.500  -0.500 1.500  ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    PORT
      LAYER ML1 ;
        POLYGON 14.800 6.200  14.800 3.200  15.800 3.200  15.800 5.200  19.800 
        5.200  19.800 12.700  20.500 12.700  20.500 14.700  19.800 14.700  
        19.800 21.100  20.000 21.100  20.000 26.500  18.600 26.500  18.600 
        21.100  18.800 21.100  18.800 14.700  18.500 14.700  18.500 12.700  
        18.800 12.700  18.800 6.200  14.800 6.200  ;
    END
  END Y
  OBS
    LAYER CNT ;
      POLYGON 17.800 3.200  17.800 4.200  18.800 4.200  18.800 3.200  17.800 
      3.200  ;
      POLYGON 18.800 23.300  18.800 24.300  19.800 24.300  19.800 23.300  
      18.800 23.300  ;
      POLYGON 18.800 21.300  18.800 22.300  19.800 22.300  19.800 21.300  
      18.800 21.300  ;
      POLYGON 18.800 25.300  18.800 26.300  19.800 26.300  19.800 25.300  
      18.800 25.300  ;
      POLYGON 6.500 14.200  6.500 15.200  7.500 15.200  7.500 14.200  6.500 
      14.200  ;
      POLYGON 9.700 29.000  9.700 30.000  10.700 30.000  10.700 29.000  9.700 
      29.000  ;
      POLYGON 16.500 7.700  16.500 8.700  17.500 8.700  17.500 7.700  16.500 
      7.700  ;
      POLYGON 13.800 14.200  13.800 15.200  14.800 15.200  14.800 14.200  
      13.800 14.200  ;
      POLYGON 3.500 10.200  3.500 11.200  4.500 11.200  4.500 10.200  3.500 
      10.200  ;
      POLYGON 10.800 10.200  10.800 11.200  11.800 11.200  11.800 10.200  
      10.800 10.200  ;
      POLYGON 9.700 0.000  9.700 1.000  10.700 1.000  10.700 0.000  9.700 
      0.000  ;
      POLYGON 15.800 23.300  15.800 24.300  16.800 24.300  16.800 23.300  
      15.800 23.300  ;
      POLYGON 15.800 25.300  15.800 26.300  16.800 26.300  16.800 25.300  
      15.800 25.300  ;
      POLYGON 15.800 21.300  15.800 22.300  16.800 22.300  16.800 21.300  
      15.800 21.300  ;
      POLYGON 14.800 3.200  14.800 4.200  15.800 4.200  15.800 3.200  14.800 
      3.200  ;
      POLYGON 12.800 25.300  12.800 26.300  13.800 26.300  13.800 25.300  
      12.800 25.300  ;
      POLYGON 12.800 23.300  12.800 24.300  13.800 24.300  13.800 23.300  
      12.800 23.300  ;
      POLYGON 12.800 21.300  12.800 22.300  13.800 22.300  13.800 21.300  
      12.800 21.300  ;
      POLYGON 9.800 3.200  9.800 4.200  10.800 4.200  10.800 3.200  9.800 
      3.200  ;
      POLYGON 9.800 25.300  9.800 26.300  10.800 26.300  10.800 25.300  9.800 
      25.300  ;
      POLYGON 9.800 23.300  9.800 24.300  10.800 24.300  10.800 23.300  9.800 
      23.300  ;
      POLYGON 9.800 21.300  9.800 22.300  10.800 22.300  10.800 21.300  9.800 
      21.300  ;
      POLYGON 7.300 3.200  7.300 4.200  8.300 4.200  8.300 3.200  7.300 3.200  ;
      
      POLYGON 6.300 25.300  6.300 26.300  7.300 26.300  7.300 25.300  6.300 
      25.300  ;
      POLYGON 6.300 21.300  6.300 22.300  7.300 22.300  7.300 21.300  6.300 
      21.300  ;
      POLYGON 6.300 23.300  6.300 24.300  7.300 24.300  7.300 23.300  6.300 
      23.300  ;
      POLYGON 4.300 3.200  4.300 4.200  5.300 4.200  5.300 3.200  4.300 3.200  ;
      
      POLYGON 1.300 25.300  1.300 26.300  2.300 26.300  2.300 25.300  1.300 
      25.300  ;
      POLYGON 1.300 3.200  1.300 4.200  2.300 4.200  2.300 3.200  1.300 3.200  ;
      
      POLYGON 1.300 21.300  1.300 22.300  2.300 22.300  2.300 21.300  1.300 
      21.300  ;
      POLYGON 1.300 23.300  1.300 24.300  2.300 24.300  2.300 23.300  1.300 
      23.300  ;
    LAYER FRAME ;
      POLYGON -0.500 1.500  -0.500 -0.500  21.500 -0.500  21.500 1.500  -0.500 
      1.500  ;
      POLYGON 0.000 0.000  21.000 0.000  21.000 30.000  0.000 30.000  0.000 
      0.000  ;
      RECT -0.500 28.500  21.500 30.500  ;
    LAYER ML1 ;
      RECT 9.200 -0.500  11.200 1.500  ;
      RECT 3.000 9.700  5.000 11.700  ;
      RECT 9.200 28.500  11.200 30.500  ;
      RECT 6.000 13.700  8.000 15.700  ;
      RECT 18.300 24.800  20.300 26.800  ;
      RECT 18.300 20.800  20.300 22.800  ;
      RECT 18.300 22.800  20.300 24.800  ;
      RECT 17.300 2.700  19.300 4.700  ;
      RECT 15.300 22.800  17.300 24.800  ;
      RECT 15.300 24.800  17.300 26.800  ;
      RECT 15.300 20.800  17.300 22.800  ;
      RECT 14.300 2.700  16.300 4.700  ;
      RECT 12.300 24.800  14.300 26.800  ;
      RECT 12.300 22.800  14.300 24.800  ;
      RECT 12.300 20.800  14.300 22.800  ;
      RECT 9.300 2.700  11.300 4.700  ;
      RECT 9.300 24.800  11.300 26.800  ;
      RECT 9.300 22.800  11.300 24.800  ;
      RECT 9.300 20.800  11.300 22.800  ;
      RECT 6.800 2.700  8.800 4.700  ;
      RECT 5.800 24.800  7.800 26.800  ;
      RECT 5.800 20.800  7.800 22.800  ;
      RECT 5.800 22.800  7.800 24.800  ;
      RECT 3.800 2.700  5.800 4.700  ;
      RECT 0.800 24.800  2.800 26.800  ;
      RECT 0.800 2.700  2.800 4.700  ;
      RECT 0.800 20.800  2.800 22.800  ;
      RECT 0.800 22.800  2.800 24.800  ;
      POLYGON -0.500 30.500  -0.500 28.500  6.100 28.500  6.100 21.900  7.500 
      21.900  7.500 28.500  12.600 28.500  12.600 21.900  14.000 21.900  
      14.000 28.500  21.500 28.500  21.500 30.500  -0.500 30.500  ;
      POLYGON -0.500 1.500  -0.500 -0.500  21.500 -0.500  21.500 1.500  18.800 
      1.500  18.800 4.200  17.800 4.200  17.800 1.500  10.800 1.500  10.800 
      4.200  9.800 4.200  9.800 1.500  8.300 1.500  8.300 4.200  7.300 4.200  
      7.300 1.500  2.300 1.500  2.300 4.200  1.300 4.200  1.300 1.500  -0.500 
      1.500  ;
      POLYGON 1.000 19.500  1.000 7.700  4.300 7.700  4.300 3.200  5.300 3.200 
       5.300 7.700  16.000 7.700  16.000 7.200  18.000 7.200  18.000 9.200  
      16.000 9.200  16.000 8.700  2.000 8.700  2.000 18.500  2.300 18.500  
      2.300 21.900  2.500 21.900  2.500 26.500  1.100 26.500  1.100 21.900  
      1.300 21.900  1.300 19.500  1.000 19.500  ;
      POLYGON 9.600 25.800  9.600 18.800  17.000 18.800  17.000 26.500  15.600 
      26.500  15.600 20.200  11.000 20.200  11.000 25.800  9.600 25.800  ;
      POLYGON 14.800 6.200  14.800 3.200  15.800 3.200  15.800 5.200  19.800 
      5.200  19.800 12.700  20.500 12.700  20.500 14.700  19.800 14.700  
      19.800 21.100  20.000 21.100  20.000 26.500  18.600 26.500  18.600 
      21.100  18.800 21.100  18.800 14.700  18.500 14.700  18.500 12.700  
      18.800 12.700  18.800 6.200  14.800 6.200  ;
      POLYGON 3.000 11.700  3.000 9.700  5.000 9.700  5.000 10.200  10.300 
      10.200  10.300 9.700  12.300 9.700  12.300 11.700  10.300 11.700  10.300 
      11.200  5.000 11.200  5.000 11.700  3.000 11.700  ;
      POLYGON 6.000 15.700  6.000 13.700  8.000 13.700  8.000 14.200  13.300 
      14.200  13.300 13.700  15.300 13.700  15.300 15.700  13.300 15.700  
      13.300 15.200  8.000 15.200  8.000 15.700  6.000 15.700  ;
    LAYER ML2 ;
      POLYGON 6.000 13.700  6.000 15.700  8.000 15.700  8.000 13.700  6.000 
      13.700  ;
      POLYGON 18.500 12.700  18.500 14.700  20.500 14.700  20.500 12.700  
      18.500 12.700  ;
      POLYGON 3.000 9.700  3.000 11.700  5.000 11.700  5.000 9.700  3.000 
      9.700  ;
    LAYER POL ;
      POLYGON 16.000 9.200  16.000 7.200  16.300 7.200  16.300 1.900  17.300 
      1.900  17.300 7.200  18.000 7.200  18.000 9.200  17.300 9.200  17.300 
      12.500  18.300 12.500  18.300 27.600  17.300 27.600  17.300 13.500  
      16.300 13.500  16.300 9.200  16.000 9.200  ;
      POLYGON 13.300 15.700  13.300 1.900  14.300 1.900  14.300 13.700  15.300 
      13.700  15.300 27.600  14.300 27.600  14.300 15.700  13.300 15.700  ;
      POLYGON 10.300 11.700  10.300 9.700  11.300 9.700  11.300 1.900  12.300 
      1.900  12.300 27.600  11.300 27.600  11.300 11.700  10.300 11.700  ;
      POLYGON 5.800 8.000  5.800 1.700  6.800 1.700  6.800 7.000  7.000 7.000  
      7.000 13.700  8.000 13.700  8.000 15.700  7.000 15.700  7.000 18.000  
      5.800 18.000  5.800 27.800  4.800 27.800  4.800 17.000  6.000 17.000  
      6.000 8.000  5.800 8.000  ;
      POLYGON 2.800 27.800  2.800 1.700  3.800 1.700  3.800 9.700  5.000 9.700 
       5.000 11.700  3.800 11.700  3.800 27.800  2.800 27.800  ;
    LAYER VIA1 ;
      POLYGON 6.500 14.200  6.500 15.200  7.500 15.200  7.500 14.200  6.500 
      14.200  ;
      POLYGON 19.000 13.200  19.000 14.200  20.000 14.200  20.000 13.200  
      19.000 13.200  ;
      POLYGON 3.500 10.200  3.500 11.200  4.500 11.200  4.500 10.200  3.500 
      10.200  ;
  END
END exorLEF


END LIBRARY
