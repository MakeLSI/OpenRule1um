VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;


MACRO cinv
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 11.500 BY 30.000 ;
  SYMMETRY X Y ;
  SITE unit ;
  
  PIN A
    USE SIGNAL ;
    PORT
      LAYER ML1 ;
        POLYGON 6.500 11.500  6.500 13.500  8.500 13.500  8.500 11.500  6.500 
        11.500  ;
    END
    PORT
      LAYER ML2 ;
        POLYGON 6.500 11.500  6.500 13.500  8.500 13.500  8.500 11.500  6.500 
        11.500  ;
    END
  END A
  PIN OE
    USE SIGNAL ;
    PORT
      LAYER ML1 ;
        POLYGON 1.000 14.500  1.000 16.500  3.000 16.500  3.000 14.500  1.000 
        14.500  ;
    END
    PORT
      LAYER ML2 ;
        POLYGON 1.000 14.500  1.000 16.500  3.000 16.500  3.000 14.500  1.000 
        14.500  ;
    END
  END OE
  PIN VDD
    USE POWER ;
    PORT
      LAYER ML1 ;
        RECT -0.500 28.500  12.000 30.500  ;
    END
  END VDD
  PIN VSS
    USE GROUND ;
    PORT
      LAYER ML1 ;
        RECT -0.500 -0.500  12.000 1.500  ;
    END
  END VSS
  PIN YB
    USE SIGNAL ;
    PORT
      LAYER ML2 ;
        POLYGON 9.000 7.200  9.000 9.200  11.000 9.200  11.000 7.200  9.000 
        7.200  ;
    END
    PORT
      LAYER ML1 ;
        POLYGON 9.000 7.200  9.000 9.200  11.000 9.200  11.000 7.200  9.000 
        7.200  ;
    END
    PORT
      LAYER ML1 ;
        WIDTH 1.000  ;
        PATH 9.800 20.500 9.800 18.000 10.000 18.000 10.000 8.200 9.800 8.200 
        9.800 3.800  ;
    END
  END YB
  OBS

    LAYER ML1 ;

      WIDTH 1.000  ;
      PATH 9.800 20.500 9.800 18.000 10.000 18.000 10.000 8.200 9.800 8.200 
      9.800 3.800  ;
      WIDTH 1.400  ;
      PATH 9.800 21.300 9.800 24.500  ;

      WIDTH 1.400  ;
      PATH 4.800 21.300 4.800 28.500  ;
      WIDTH 1.000  ;
      PATH 4.800 1.000 4.800 3.800  ;
      WIDTH 1.400  ;
      PATH 1.800 21.300 1.800 24.500  ;
      WIDTH 1.000  ;
      PATH 1.800 24.500 1.800 18.000 5.000 18.000 5.000 8.000 1.800 8.000 
      1.800 3.800  ;

    VIA 1.800 22.500  dcont ;
    VIA 1.800 20.500  dcont ;
    VIA 1.800 3.800  dcont ;
    VIA 1.800 24.500  dcont ;
    VIA 4.800 22.500  dcont ;
    VIA 4.800 20.500  dcont ;
    VIA 4.800 24.500  dcont ;
    VIA 4.800 3.800  dcont ;
    VIA 9.800 3.800  dcont ;
    VIA 9.800 20.500  dcont ;
    VIA 9.800 22.500  dcont ;
    VIA 9.800 24.500  dcont ;
    VIA 7.000 29.500  nsubcont ;
    VIA 7.500 12.500  pcont ;
    VIA 5.800 15.500  pcont ;
    VIA 2.000 15.500  pcont ;
    VIA 6.000 0.500  psubcont ;
  END
END cinv

MACRO dcont
  CLASS CORE ;
  OBS
    LAYER ML1 ;
      RECT -1.000 -1.000  1.000 1.000  ;
  END
END dcont

MACRO nsubcont
  CLASS CORE ;
  OBS
    LAYER ML1 ;
      RECT -1.000 -1.000  1.000 1.000  ;
  END
END nsubcont

MACRO pcont
  CLASS CORE ;
  OBS
    LAYER ML1 ;
      RECT -1.000 -1.000  1.000 1.000  ;
  END
END pcont

MACRO psubcont
  CLASS CORE ;
  OBS
    LAYER ML1 ;
      RECT -1.000 -1.000  1.000 1.000  ;
  END
END psubcont


END LIBRARY
