VERSION 5.3 ;

NAMESCASESENSITIVE ON ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS











MACRO na212LEF
  CLASS BLOCK ;
  PIN A0
    DIRECTION INPUT ;
    PORT
      LAYER POL ;
        POLYGON 1.000 16.500  1.000 14.500  2.000 14.500  2.000 9.500  2.800 
        9.500  2.800 3.500  3.800 3.500  3.800 10.500  3.000 10.500  3.000 
        17.100  4.800 17.100  4.800 26.500  3.800 26.500  3.800 18.100  2.000 
        18.100  2.000 16.500  1.000 16.500  ;
    END
    PORT
      LAYER ML1 ;
        POLYGON 1.000 14.500  1.000 16.500  3.000 16.500  3.000 14.500  1.000 
        14.500  ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER POL ;
        POLYGON 4.000 13.500  4.000 11.500  5.000 11.500  5.000 9.500  5.800 
        9.500  5.800 3.500  6.800 3.500  6.800 10.500  6.000 10.500  6.000 
        15.000  6.800 15.000  6.800 26.500  5.800 26.500  5.800 16.000  5.000 
        16.000  5.000 13.500  4.000 13.500  ;
    END
    PORT
      LAYER ML1 ;
        POLYGON 4.000 11.500  4.000 13.500  6.000 13.500  6.000 11.500  4.000 
        11.500  ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    PORT
      LAYER POL ;
        POLYGON 7.000 14.000  7.000 12.000  8.800 12.000  8.800 3.500  9.800 
        3.500  9.800 13.400  9.000 13.400  9.000 17.500  9.800 17.500  9.800 
        26.500  8.800 26.500  8.800 18.500  8.000 18.500  8.000 14.000  7.000 
        14.000  ;
    END
    PORT
      LAYER ML1 ;
        POLYGON 7.000 12.000  7.000 14.000  9.000 14.000  9.000 12.000  7.000 
        12.000  ;
    END
  END B0
  PIN VDD
    DIRECTION INOUT ;
    PORT
      LAYER ML1 ;
        POLYGON -0.500 30.500  -0.500 28.500  2.100 28.500  2.100 20.600  
        3.500 20.600  3.500 28.500  10.100 28.500  10.100 20.600  11.500 
        20.600  11.500 28.500  13.000 28.500  13.000 30.500  -0.500 30.500  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    PORT
      LAYER ML1 ;
        POLYGON -0.500 1.500  -0.500 -0.500  13.000 -0.500  13.000 1.500  
        5.300 1.500  5.300 6.000  4.300 6.000  4.300 1.500  -0.500 1.500  ;
    END
  END VSS
  PIN YB
    DIRECTION OUTPUT ;
    PORT
      LAYER ML1 ;
        POLYGON 7.100 25.200  7.100 20.600  7.300 20.600  7.300 17.500  10.000 
        17.500  10.000 7.500  10.300 7.500  10.300 5.000  11.300 5.000  11.300 
        8.500  12.000 8.500  12.000 10.500  11.000 10.500  11.000 18.500  
        8.300 18.500  8.300 20.600  8.500 20.600  8.500 25.200  7.100 25.200  ;
    END
  END YB
  OBS
    LAYER CNT ;
      POLYGON 7.300 20.000  7.300 21.000  8.300 21.000  8.300 20.000  7.300 
      20.000  ;
      POLYGON 7.300 5.000  7.300 6.000  8.300 6.000  8.300 5.000  7.300 5.000  ;
      
      POLYGON 10.300 5.000  10.300 6.000  11.300 6.000  11.300 5.000  10.300 
      5.000  ;
      POLYGON 10.300 20.000  10.300 21.000  11.300 21.000  11.300 20.000  
      10.300 20.000  ;
      POLYGON 10.300 22.000  10.300 23.000  11.300 23.000  11.300 22.000  
      10.300 22.000  ;
      POLYGON 10.300 24.000  10.300 25.000  11.300 25.000  11.300 24.000  
      10.300 24.000  ;
      POLYGON 7.500 12.500  7.500 13.500  8.500 13.500  8.500 12.500  7.500 
      12.500  ;
      POLYGON 7.700 29.000  7.700 30.000  8.700 30.000  8.700 29.000  7.700 
      29.000  ;
      POLYGON 4.500 12.000  4.500 13.000  5.500 13.000  5.500 12.000  4.500 
      12.000  ;
      POLYGON 1.500 15.000  1.500 16.000  2.500 16.000  2.500 15.000  1.500 
      15.000  ;
      POLYGON 6.000 0.000  6.000 1.000  7.000 1.000  7.000 0.000  6.000 0.000  ;
      
      POLYGON 7.300 22.000  7.300 23.000  8.300 23.000  8.300 22.000  7.300 
      22.000  ;
      POLYGON 7.300 24.000  7.300 25.000  8.300 25.000  8.300 24.000  7.300 
      24.000  ;
      POLYGON 4.300 5.000  4.300 6.000  5.300 6.000  5.300 5.000  4.300 5.000  ;
      
      POLYGON 2.300 24.000  2.300 25.000  3.300 25.000  3.300 24.000  2.300 
      24.000  ;
      POLYGON 2.300 20.000  2.300 21.000  3.300 21.000  3.300 20.000  2.300 
      20.000  ;
      POLYGON 2.300 22.000  2.300 23.000  3.300 23.000  3.300 22.000  2.300 
      22.000  ;
      POLYGON 1.300 5.000  1.300 6.000  2.300 6.000  2.300 5.000  1.300 5.000  ;
      
    LAYER FRAME ;
      RECT -0.500 28.500  13.000 30.500  ;
      RECT -0.500 -0.500  13.000 1.500  ;
      POLYGON 0.000 0.000  12.500 0.000  12.500 30.000  0.000 30.000  0.000 
      0.000  ;
    LAYER ML1 ;
      POLYGON 4.000 11.500  4.000 13.500  6.000 13.500  6.000 11.500  4.000 
      11.500  ;
      POLYGON 1.000 14.500  1.000 16.500  3.000 16.500  3.000 14.500  1.000 
      14.500  ;
      RECT 5.500 -0.500  7.500 1.500  ;
      POLYGON 7.000 12.000  7.000 14.000  9.000 14.000  9.000 12.000  7.000 
      12.000  ;
      RECT 1.000 14.500  3.000 16.500  ;
      RECT 4.000 11.500  6.000 13.500  ;
      RECT 7.200 28.500  9.200 30.500  ;
      RECT 7.000 12.000  9.000 14.000  ;
      RECT 9.800 23.500  11.800 25.500  ;
      RECT 9.800 21.500  11.800 23.500  ;
      RECT 9.800 19.500  11.800 21.500  ;
      RECT 9.800 4.500  11.800 6.500  ;
      RECT 6.800 4.500  8.800 6.500  ;
      RECT 6.800 19.500  8.800 21.500  ;
      RECT 6.800 21.500  8.800 23.500  ;
      RECT 6.800 23.500  8.800 25.500  ;
      RECT 3.800 4.500  5.800 6.500  ;
      RECT 1.800 23.500  3.800 25.500  ;
      RECT 1.800 19.500  3.800 21.500  ;
      RECT 1.800 21.500  3.800 23.500  ;
      RECT 0.800 4.500  2.800 6.500  ;
      POLYGON -0.500 30.500  -0.500 28.500  2.100 28.500  2.100 20.600  3.500 
      20.600  3.500 28.500  10.100 28.500  10.100 20.600  11.500 20.600  
      11.500 28.500  13.000 28.500  13.000 30.500  -0.500 30.500  ;
      POLYGON 7.100 25.200  7.100 20.600  7.300 20.600  7.300 17.500  10.000 
      17.500  10.000 7.500  10.300 7.500  10.300 5.000  11.300 5.000  11.300 
      8.500  12.000 8.500  12.000 10.500  11.000 10.500  11.000 18.500  8.300 
      18.500  8.300 20.600  8.500 20.600  8.500 25.200  7.100 25.200  ;
      POLYGON 1.300 8.500  1.300 5.000  2.300 5.000  2.300 7.500  7.300 7.500  
      7.300 5.000  8.300 5.000  8.300 8.500  1.300 8.500  ;
      POLYGON -0.500 1.500  -0.500 -0.500  13.000 -0.500  13.000 1.500  5.300 
      1.500  5.300 6.000  4.300 6.000  4.300 1.500  -0.500 1.500  ;
    LAYER ML2 ;
      POLYGON 10.000 10.500  10.000 8.500  12.000 8.500  12.000 10.500  10.000 
      10.500  ;
      POLYGON 7.000 12.000  7.000 14.000  9.000 14.000  9.000 12.000  7.000 
      12.000  ;
      POLYGON 4.000 11.500  4.000 13.500  6.000 13.500  6.000 11.500  4.000 
      11.500  ;
      POLYGON 1.000 14.500  1.000 16.500  3.000 16.500  3.000 14.500  1.000 
      14.500  ;
    LAYER POL ;
      POLYGON 7.000 14.000  7.000 12.000  8.800 12.000  8.800 3.500  9.800 
      3.500  9.800 13.400  9.000 13.400  9.000 17.500  9.800 17.500  9.800 
      26.500  8.800 26.500  8.800 18.500  8.000 18.500  8.000 14.000  7.000 
      14.000  ;
      POLYGON 4.000 13.500  4.000 11.500  5.000 11.500  5.000 9.500  5.800 
      9.500  5.800 3.500  6.800 3.500  6.800 10.500  6.000 10.500  6.000 
      15.000  6.800 15.000  6.800 26.500  5.800 26.500  5.800 16.000  5.000 
      16.000  5.000 13.500  4.000 13.500  ;
      POLYGON 1.000 16.500  1.000 14.500  2.000 14.500  2.000 9.500  2.800 
      9.500  2.800 3.500  3.800 3.500  3.800 10.500  3.000 10.500  3.000 
      17.100  4.800 17.100  4.800 26.500  3.800 26.500  3.800 18.100  2.000 
      18.100  2.000 16.500  1.000 16.500  ;
    LAYER VIA1 ;
      POLYGON 7.500 12.500  7.500 13.500  8.500 13.500  8.500 12.500  7.500 
      12.500  ;
      POLYGON 4.500 12.000  4.500 13.000  5.500 13.000  5.500 12.000  4.500 
      12.000  ;
      POLYGON 10.500 9.000  10.500 10.000  11.500 10.000  11.500 9.000  10.500 
      9.000  ;
      POLYGON 1.500 15.000  1.500 16.000  2.500 16.000  2.500 15.000  1.500 
      15.000  ;
  END
END na212LEF


END LIBRARY
