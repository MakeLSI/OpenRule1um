VERSION 5.3 ;

NAMESCASESENSITIVE ON ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS











MACRO na31LEF
  CLASS BLOCK ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER POL ;
        POLYGON 1.000 16.500  1.000 14.500  2.000 14.500  2.000 6.000  2.800 
        6.000  2.800 1.700  3.800 1.700  3.800 7.000  3.000 7.000  3.000 
        15.000  3.800 15.000  3.800 26.500  2.800 26.500  2.800 16.500  1.000 
        16.500  ;
    END
    PORT
      LAYER ML1 ;
        POLYGON 1.000 14.500  1.000 16.500  3.000 16.500  3.000 14.500  1.000 
        14.500  ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER POL ;
        POLYGON 4.000 13.500  4.000 11.500  4.800 11.500  4.800 1.700  5.800 
        1.700  5.800 11.500  6.000 11.500  6.000 15.000  6.800 15.000  6.800 
        26.500  5.800 26.500  5.800 16.000  5.000 16.000  5.000 13.500  4.000 
        13.500  ;
    END
    PORT
      LAYER ML1 ;
        POLYGON 4.000 11.500  4.000 13.500  6.000 13.500  6.000 11.500  4.000 
        11.500  ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER POL ;
        POLYGON 6.800 9.000  6.800 1.700  7.800 1.700  7.800 8.000  9.800 
        8.000  9.800 26.500  8.800 26.500  8.800 9.000  6.800 9.000  ;
    END
    PORT
      LAYER ML1 ;
        POLYGON 7.000 10.000  7.000 8.000  9.000 8.000  9.000 10.000  7.000 
        10.000  ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    PORT
      LAYER ML1 ;
        POLYGON -0.500 30.500  -0.500 28.500  1.100 28.500  1.100 20.600  
        2.500 20.600  2.500 28.500  7.100 28.500  7.100 20.600  8.500 20.600  
        8.500 28.500  13.000 28.500  13.000 30.500  -0.500 30.500  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    PORT
      LAYER ML1 ;
        POLYGON -0.500 1.500  -0.500 -0.500  13.000 -0.500  13.000 1.500  
        2.300 1.500  2.300 4.200  1.300 4.200  1.300 1.500  -0.500 1.500  ;
    END
  END VSS
  PIN YB
    DIRECTION OUTPUT ;
    PORT
      LAYER ML1 ;
        POLYGON 8.300 7.000  8.300 3.200  9.300 3.200  9.300 6.000  11.300 
        6.000  11.300 12.000  12.000 12.000  12.000 14.000  11.300 14.000  
        11.300 20.600  11.500 20.600  11.500 25.200  10.100 25.200  10.100 
        20.600  10.300 20.600  10.300 18.500  5.300 18.500  5.300 20.600  
        5.500 20.600  5.500 25.200  4.100 25.200  4.100 20.600  4.300 20.600  
        4.300 17.500  10.300 17.500  10.300 14.000  10.000 14.000  10.000 
        12.000  10.300 12.000  10.300 7.000  8.300 7.000  ;
    END
  END YB
  OBS
    LAYER CNT ;
      POLYGON 7.300 22.000  7.300 23.000  8.300 23.000  8.300 22.000  7.300 
      22.000  ;
      POLYGON 7.300 20.000  7.300 21.000  8.300 21.000  8.300 20.000  7.300 
      20.000  ;
      POLYGON 8.300 3.200  8.300 4.200  9.300 4.200  9.300 3.200  8.300 3.200  ;
      
      POLYGON 10.300 24.000  10.300 25.000  11.300 25.000  11.300 24.000  
      10.300 24.000  ;
      POLYGON 10.300 22.000  10.300 23.000  11.300 23.000  11.300 22.000  
      10.300 22.000  ;
      POLYGON 10.300 20.000  10.300 21.000  11.300 21.000  11.300 20.000  
      10.300 20.000  ;
      POLYGON 7.500 8.500  7.500 9.500  8.500 9.500  8.500 8.500  7.500 8.500  ;
      
      POLYGON 5.000 29.000  5.000 30.000  6.000 30.000  6.000 29.000  5.000 
      29.000  ;
      POLYGON 4.500 12.000  4.500 13.000  5.500 13.000  5.500 12.000  4.500 
      12.000  ;
      POLYGON 1.500 15.000  1.500 16.000  2.500 16.000  2.500 15.000  1.500 
      15.000  ;
      POLYGON 4.500 0.000  4.500 1.000  5.500 1.000  5.500 0.000  4.500 0.000  ;
      
      POLYGON 7.300 24.000  7.300 25.000  8.300 25.000  8.300 24.000  7.300 
      24.000  ;
      POLYGON 4.300 24.000  4.300 25.000  5.300 25.000  5.300 24.000  4.300 
      24.000  ;
      POLYGON 4.300 20.000  4.300 21.000  5.300 21.000  5.300 20.000  4.300 
      20.000  ;
      POLYGON 4.300 22.000  4.300 23.000  5.300 23.000  5.300 22.000  4.300 
      22.000  ;
      POLYGON 1.300 24.000  1.300 25.000  2.300 25.000  2.300 24.000  1.300 
      24.000  ;
      POLYGON 1.300 3.200  1.300 4.200  2.300 4.200  2.300 3.200  1.300 3.200  ;
      
      POLYGON 1.300 20.000  1.300 21.000  2.300 21.000  2.300 20.000  1.300 
      20.000  ;
      POLYGON 1.300 22.000  1.300 23.000  2.300 23.000  2.300 22.000  1.300 
      22.000  ;
    LAYER FRAME ;
      RECT -0.500 28.500  13.000 30.500  ;
      RECT -0.500 -0.500  13.000 1.500  ;
      POLYGON 0.000 0.000  12.500 0.000  12.500 30.000  0.000 30.000  0.000 
      0.000  ;
    LAYER ML1 ;
      POLYGON 1.000 14.500  1.000 16.500  3.000 16.500  3.000 14.500  1.000 
      14.500  ;
      POLYGON 4.000 11.500  4.000 13.500  6.000 13.500  6.000 11.500  4.000 
      11.500  ;
      RECT 4.000 -0.500  6.000 1.500  ;
      RECT 1.000 14.500  3.000 16.500  ;
      RECT 4.000 11.500  6.000 13.500  ;
      RECT 4.500 28.500  6.500 30.500  ;
      RECT 7.000 8.000  9.000 10.000  ;
      RECT 9.800 19.500  11.800 21.500  ;
      RECT 9.800 21.500  11.800 23.500  ;
      RECT 9.800 23.500  11.800 25.500  ;
      RECT 7.800 2.700  9.800 4.700  ;
      RECT 6.800 19.500  8.800 21.500  ;
      RECT 6.800 21.500  8.800 23.500  ;
      RECT 6.800 23.500  8.800 25.500  ;
      RECT 3.800 23.500  5.800 25.500  ;
      RECT 3.800 19.500  5.800 21.500  ;
      RECT 3.800 21.500  5.800 23.500  ;
      RECT 0.800 23.500  2.800 25.500  ;
      RECT 0.800 2.700  2.800 4.700  ;
      RECT 0.800 19.500  2.800 21.500  ;
      RECT 0.800 21.500  2.800 23.500  ;
      POLYGON -0.500 30.500  -0.500 28.500  1.100 28.500  1.100 20.600  2.500 
      20.600  2.500 28.500  7.100 28.500  7.100 20.600  8.500 20.600  8.500 
      28.500  13.000 28.500  13.000 30.500  -0.500 30.500  ;
      POLYGON -0.500 1.500  -0.500 -0.500  13.000 -0.500  13.000 1.500  2.300 
      1.500  2.300 4.200  1.300 4.200  1.300 1.500  -0.500 1.500  ;
      POLYGON 8.300 7.000  8.300 3.200  9.300 3.200  9.300 6.000  11.300 6.000 
       11.300 12.000  12.000 12.000  12.000 14.000  11.300 14.000  11.300 
      20.600  11.500 20.600  11.500 25.200  10.100 25.200  10.100 20.600  
      10.300 20.600  10.300 18.500  5.300 18.500  5.300 20.600  5.500 20.600  
      5.500 25.200  4.100 25.200  4.100 20.600  4.300 20.600  4.300 17.500  
      10.300 17.500  10.300 14.000  10.000 14.000  10.000 12.000  10.300 
      12.000  10.300 7.000  8.300 7.000  ;
      POLYGON 7.000 10.000  7.000 8.000  9.000 8.000  9.000 10.000  7.000 
      10.000  ;
    LAYER ML2 ;
      POLYGON 10.000 14.000  10.000 12.000  12.000 12.000  12.000 14.000  
      10.000 14.000  ;
      POLYGON 7.000 8.000  7.000 10.000  9.000 10.000  9.000 8.000  7.000 
      8.000  ;
      POLYGON 4.000 11.500  4.000 13.500  6.000 13.500  6.000 11.500  4.000 
      11.500  ;
      POLYGON 1.000 14.500  1.000 16.500  3.000 16.500  3.000 14.500  1.000 
      14.500  ;
    LAYER POL ;
      POLYGON 6.800 9.000  6.800 1.700  7.800 1.700  7.800 8.000  9.800 8.000  
      9.800 26.500  8.800 26.500  8.800 9.000  6.800 9.000  ;
      POLYGON 4.000 13.500  4.000 11.500  4.800 11.500  4.800 1.700  5.800 
      1.700  5.800 11.500  6.000 11.500  6.000 15.000  6.800 15.000  6.800 
      26.500  5.800 26.500  5.800 16.000  5.000 16.000  5.000 13.500  4.000 
      13.500  ;
      POLYGON 1.000 16.500  1.000 14.500  2.000 14.500  2.000 6.000  2.800 
      6.000  2.800 1.700  3.800 1.700  3.800 7.000  3.000 7.000  3.000 15.000  
      3.800 15.000  3.800 26.500  2.800 26.500  2.800 16.500  1.000 16.500  ;
      POLYGON 7.000 8.000  7.000 10.000  9.000 10.000  9.000 8.000  7.000 
      8.000  ;
    LAYER VIA1 ;
      POLYGON 7.500 8.500  7.500 9.500  8.500 9.500  8.500 8.500  7.500 8.500  ;
      
      POLYGON 4.500 12.000  4.500 13.000  5.500 13.000  5.500 12.000  4.500 
      12.000  ;
      POLYGON 10.500 12.500  10.500 13.500  11.500 13.500  11.500 12.500  
      10.500 12.500  ;
      POLYGON 1.500 15.000  1.500 16.000  2.500 16.000  2.500 15.000  1.500 
      15.000  ;
  END
END na31LEF


END LIBRARY
