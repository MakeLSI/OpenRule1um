VERSION 5.3 ;

NAMESCASESENSITIVE ON ;

BUSBITCHARS "[]" ;

DIVIDERCHAR "/" ;

LAYER Via
 TYPE CUT ;
 WIDTH 0.600 ;
 SPACING 0.600  ;
END Via

LAYER Via2
 TYPE CUT ;
 WIDTH 0.600 ;
 SPACING 0.600  ;
END Via2

LAYER M1
 TYPE ROUTING ;
 WIDTH 0.800 ;
 PITCH 0.050 ;
 OFFSET 0.000 ;
 SPACING 0.800 ;
 RESISTANCE RPERSQ 0.000000e+000 ;
 CAPACITANCE CPERSQDIST 0.000000e+000 ;
 EDGECAPACITANCE 0.000000e+000 ;
 ANTENNAAREAFACTOR 0.000000 ;
 ANTENNALENGTHFACTOR 0.000000 ;
END M1

LAYER M2
 TYPE ROUTING ;
 WIDTH 0.800 ;
 PITCH 0.050 ;
 OFFSET 0.000 ;
 SPACING 0.800 ;
 RESISTANCE RPERSQ 0.000000e+000 ;
 CAPACITANCE CPERSQDIST 0.000000e+000 ;
 EDGECAPACITANCE 0.000000e+000 ;
 ANTENNAAREAFACTOR 0.000000 ;
 ANTENNALENGTHFACTOR 0.000000 ;
END M2

LAYER M3
 TYPE ROUTING ;
 WIDTH 0.800 ;
 PITCH 0.050 ;
 OFFSET 0.000 ;
 SPACING 0.800 ;
 RESISTANCE RPERSQ 0.000000e+000 ;
 CAPACITANCE CPERSQDIST 0.000000e+000 ;
 EDGECAPACITANCE 0.000000e+000 ;
 ANTENNAAREAFACTOR 0.000000 ;
 ANTENNALENGTHFACTOR 0.000000 ;
END M3

LAYER Poly
 TYPE ROUTING ;
 WIDTH 0.600 ;
 PITCH 0.050 ;
 OFFSET 0.000 ;
 SPACING 0.600 ;
 RESISTANCE RPERSQ 0.000000e+000 ;
 CAPACITANCE CPERSQDIST 0.000000e+000 ;
 EDGECAPACITANCE 0.000000e+000 ;
 ANTENNAAREAFACTOR 0.000000 ;
 ANTENNALENGTHFACTOR 0.000000 ;
END Poly

LAYER Cont
 TYPE CUT ;
 WIDTH 0.600 ;
 SPACING 0.600  ;
END Cont

LAYER Diff
 TYPE ROUTING ;
 WIDTH 0.800 ;
 PITCH 0.050 ;
 OFFSET 0.000 ;
 SPACING 1.200 ;
 RESISTANCE RPERSQ 0.000000e+000 ;
 CAPACITANCE CPERSQDIST 0.000000e+000 ;
 EDGECAPACITANCE 0.000000e+000 ;
 ANTENNAAREAFACTOR 0.000000 ;
 ANTENNALENGTHFACTOR 0.000000 ;
END Diff



VIARULE PCNT
 LAYER Poly ;
 LAYER M1 ;
 VIA PCNT ;
END PCNT

VIARULE VIA12
 LAYER M1 ;
 LAYER M2 ;
 VIA VIA12 ;
END VIA12

VIARULE VIA23
 LAYER M2 ;
 LAYER M3 ;
 VIA VIA23 ;
END VIA23

VIARULE TANSHIT
 LAYER Poly ;
 LAYER M1 ;
 VIA TANSHIT ;
END TANSHIT

VIARULE POLCNT_VIAGEN_
 LAYER Poly ;
  OVERHANG 0.400 ;
 LAYER M1 ;
  OVERHANG 0.300 ;
END POLCNT_VIAGEN_

VIARULE VIA12_VIAGEN_
 LAYER M1 ;
  OVERHANG 0.400 ;
 LAYER M2 ;
  OVERHANG 4.000 ;
 VIA R ;
END VIA12_VIAGEN_










SPACING
 SAMENET FRAME Diff 0.600 ;
 SAMENET FRAME M1 0.400 ;
 SAMENET FRAME M2 0.400 ;
END SPACING





END LIBRARY
