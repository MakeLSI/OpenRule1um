VERSION 5.3 ;

NAMESCASESENSITIVE ON ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS











MACRO dff1m2LEF
  CLASS BLOCK ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER POL ;
        POLYGON 2.800 27.800  2.800 1.700  3.800 1.700  3.800 9.000  5.300 
        9.000  5.300 11.000  3.800 11.000  3.800 27.800  2.800 27.800  ;
    END
    PORT
      LAYER ML1 ;
        POLYGON 3.300 9.000  3.300 11.000  5.300 11.000  5.300 9.000  3.300 
        9.000  ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER POL ;
        POLYGON 11.000 11.000  11.000 9.000  12.300 9.000  12.300 1.900  
        13.300 1.900  13.300 27.600  12.300 27.600  12.300 11.000  11.000 
        11.000  ;
    END
    PORT
      LAYER ML1 ;
        POLYGON 11.000 9.000  11.000 11.000  13.000 11.000  13.000 9.000  
        11.000 9.000  ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER ML1 ;
        POLYGON 49.500 12.500  49.500 10.500  50.300 10.500  50.300 2.700  
        51.300 2.700  51.300 10.500  51.500 10.500  51.500 12.500  51.300 
        12.500  51.300 26.500  50.300 26.500  50.300 12.500  49.500 12.500  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    PORT
      LAYER ML1 ;
        POLYGON -0.500 30.500  -0.500 28.500  4.100 28.500  4.100 21.900  
        5.500 21.900  5.500 28.500  10.600 28.500  10.600 21.900  12.000 
        21.900  12.000 28.500  20.600 28.500  20.600 21.900  22.000 21.900  
        22.000 28.500  27.100 28.500  27.100 21.100  28.500 21.100  28.500 
        28.500  37.100 28.500  37.100 21.900  38.500 21.900  38.500 28.500  
        46.600 28.500  46.600 21.900  48.000 21.900  48.000 28.500  52.500 
        28.500  52.500 30.500  -0.500 30.500  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    PORT
      LAYER ML1 ;
        POLYGON -0.500 1.500  -0.500 -0.500  52.500 -0.500  52.500 1.500  
        48.000 1.500  48.000 4.400  46.600 4.400  46.600 1.500  38.500 1.500  
        38.500 4.400  37.100 4.400  37.100 1.500  28.500 1.500  28.500 4.400  
        27.100 4.400  27.100 1.500  22.000 1.500  22.000 4.400  20.600 4.400  
        20.600 1.500  12.000 1.500  12.000 4.400  10.600 4.400  10.600 1.500  
        5.500 1.500  5.500 4.400  4.100 4.400  4.100 1.500  -0.500 1.500  ;
    END
  END VSS
  OBS
    LAYER CNT ;
      POLYGON 33.300 13.200  33.300 14.200  34.300 14.200  34.300 13.200  
      33.300 13.200  ;
      POLYGON 36.300 13.500  36.300 14.500  37.300 14.500  37.300 13.500  
      36.300 13.500  ;
      POLYGON 38.300 18.200  38.300 19.200  39.300 19.200  39.300 18.200  
      38.300 18.200  ;
      POLYGON 38.300 6.200  38.300 7.200  39.300 7.200  39.300 6.200  38.300 
      6.200  ;
      POLYGON 44.800 8.200  44.800 9.200  45.800 9.200  45.800 8.200  44.800 
      8.200  ;
      POLYGON 44.800 16.700  44.800 17.700  45.800 17.700  45.800 16.700  
      44.800 16.700  ;
      POLYGON 47.800 6.200  47.800 7.200  48.800 7.200  48.800 6.200  47.800 
      6.200  ;
      POLYGON 47.800 18.400  47.800 19.400  48.800 19.400  48.800 18.400  
      47.800 18.400  ;
      POLYGON 45.500 0.000  45.500 1.000  46.500 1.000  46.500 0.000  45.500 
      0.000  ;
      POLYGON 27.200 0.000  27.200 1.000  28.200 1.000  28.200 0.000  27.200 
      0.000  ;
      POLYGON 9.700 0.000  9.700 1.000  10.700 1.000  10.700 0.000  9.700 
      0.000  ;
      POLYGON 31.300 16.200  31.300 17.200  32.300 17.200  32.300 16.200  
      31.300 16.200  ;
      POLYGON 28.300 12.500  28.300 13.500  29.300 13.500  29.300 12.500  
      28.300 12.500  ;
      POLYGON 24.800 18.200  24.800 19.200  25.800 19.200  25.800 18.200  
      24.800 18.200  ;
      POLYGON 24.300 6.200  24.300 7.200  25.300 7.200  25.300 6.200  24.300 
      6.200  ;
      POLYGON 21.800 9.500  21.800 10.500  22.800 10.500  22.800 9.500  21.800 
      9.500  ;
      POLYGON 21.800 18.200  21.800 19.200  22.800 19.200  22.800 18.200  
      21.800 18.200  ;
      POLYGON 19.800 6.200  19.800 7.200  20.800 7.200  20.800 6.200  19.800 
      6.200  ;
      POLYGON 16.800 15.500  16.800 16.500  17.800 16.500  17.800 15.500  
      16.800 15.500  ;
      POLYGON 14.800 12.500  14.800 13.500  15.800 13.500  15.800 12.500  
      14.800 12.500  ;
      POLYGON 14.300 6.200  14.300 7.200  15.300 7.200  15.300 6.200  14.300 
      6.200  ;
      POLYGON 11.500 9.500  11.500 10.500  12.500 10.500  12.500 9.500  11.500 
      9.500  ;
      POLYGON 9.800 12.500  9.800 13.500  10.800 13.500  10.800 12.500  9.800 
      12.500  ;
      POLYGON 5.300 6.200  5.300 7.200  6.300 7.200  6.300 6.200  5.300 6.200  ;
      
      POLYGON 5.300 18.300  5.300 19.300  6.300 19.300  6.300 18.300  5.300 
      18.300  ;
      POLYGON 4.800 12.500  4.800 13.500  5.800 13.500  5.800 12.500  4.800 
      12.500  ;
      POLYGON 3.800 9.500  3.800 10.500  4.800 10.500  4.800 9.500  3.800 
      9.500  ;
      POLYGON 9.700 29.000  9.700 30.000  10.700 30.000  10.700 29.000  9.700 
      29.000  ;
      POLYGON 27.200 29.000  27.200 30.000  28.200 30.000  28.200 29.000  
      27.200 29.000  ;
      POLYGON 45.500 29.000  45.500 30.000  46.500 30.000  46.500 29.000  
      45.500 29.000  ;
      POLYGON 49.800 25.300  49.800 26.300  50.800 26.300  50.800 25.300  
      49.800 25.300  ;
      POLYGON 49.800 23.300  49.800 24.300  50.800 24.300  50.800 23.300  
      49.800 23.300  ;
      POLYGON 49.800 21.300  49.800 22.300  50.800 22.300  50.800 21.300  
      49.800 21.300  ;
      POLYGON 49.800 3.200  49.800 4.200  50.800 4.200  50.800 3.200  49.800 
      3.200  ;
      POLYGON 46.800 25.300  46.800 26.300  47.800 26.300  47.800 25.300  
      46.800 25.300  ;
      POLYGON 46.800 23.300  46.800 24.300  47.800 24.300  47.800 23.300  
      46.800 23.300  ;
      POLYGON 46.800 21.300  46.800 22.300  47.800 22.300  47.800 21.300  
      46.800 21.300  ;
      POLYGON 46.800 3.200  46.800 4.200  47.800 4.200  47.800 3.200  46.800 
      3.200  ;
      POLYGON 43.800 25.300  43.800 26.300  44.800 26.300  44.800 25.300  
      43.800 25.300  ;
      POLYGON 43.800 23.300  43.800 24.300  44.800 24.300  44.800 23.300  
      43.800 23.300  ;
      POLYGON 43.800 21.300  43.800 22.300  44.800 22.300  44.800 21.300  
      43.800 21.300  ;
      POLYGON 43.800 3.200  43.800 4.200  44.800 4.200  44.800 3.200  43.800 
      3.200  ;
      POLYGON 40.300 3.200  40.300 4.200  41.300 4.200  41.300 3.200  40.300 
      3.200  ;
      POLYGON 40.300 25.300  40.300 26.300  41.300 26.300  41.300 25.300  
      40.300 25.300  ;
      POLYGON 40.300 23.300  40.300 24.300  41.300 24.300  41.300 23.300  
      40.300 23.300  ;
      POLYGON 40.300 21.300  40.300 22.300  41.300 22.300  41.300 21.300  
      40.300 21.300  ;
      POLYGON 37.300 3.200  37.300 4.200  38.300 4.200  38.300 3.200  37.300 
      3.200  ;
      POLYGON 37.300 25.300  37.300 26.300  38.300 26.300  38.300 25.300  
      37.300 25.300  ;
      POLYGON 37.300 23.300  37.300 24.300  38.300 24.300  38.300 23.300  
      37.300 23.300  ;
      POLYGON 37.300 21.300  37.300 22.300  38.300 22.300  38.300 21.300  
      37.300 21.300  ;
      POLYGON 32.300 3.200  32.300 4.200  33.300 4.200  33.300 3.200  32.300 
      3.200  ;
      POLYGON 32.300 25.300  32.300 26.300  33.300 26.300  33.300 25.300  
      32.300 25.300  ;
      POLYGON 32.300 23.300  32.300 24.300  33.300 24.300  33.300 23.300  
      32.300 23.300  ;
      POLYGON 32.300 21.300  32.300 22.300  33.300 22.300  33.300 21.300  
      32.300 21.300  ;
      POLYGON 27.300 3.200  27.300 4.200  28.300 4.200  28.300 3.200  27.300 
      3.200  ;
      POLYGON 27.300 23.300  27.300 24.300  28.300 24.300  28.300 23.300  
      27.300 23.300  ;
      POLYGON 27.300 25.300  27.300 26.300  28.300 26.300  28.300 25.300  
      27.300 25.300  ;
      POLYGON 23.800 3.200  23.800 4.200  24.800 4.200  24.800 3.200  23.800 
      3.200  ;
      POLYGON 23.800 25.300  23.800 26.300  24.800 26.300  24.800 25.300  
      23.800 25.300  ;
      POLYGON 23.800 23.300  23.800 24.300  24.800 24.300  24.800 23.300  
      23.800 23.300  ;
      POLYGON 20.800 3.200  20.800 4.200  21.800 4.200  21.800 3.200  20.800 
      3.200  ;
      POLYGON 20.800 25.300  20.800 26.300  21.800 26.300  21.800 25.300  
      20.800 25.300  ;
      POLYGON 20.800 23.300  20.800 24.300  21.800 24.300  21.800 23.300  
      20.800 23.300  ;
      POLYGON 20.800 21.300  20.800 22.300  21.800 22.300  21.800 21.300  
      20.800 21.300  ;
      POLYGON 15.800 3.200  15.800 4.200  16.800 4.200  16.800 3.200  15.800 
      3.200  ;
      POLYGON 15.800 23.300  15.800 24.300  16.800 24.300  16.800 23.300  
      15.800 23.300  ;
      POLYGON 15.800 25.300  15.800 26.300  16.800 26.300  16.800 25.300  
      15.800 25.300  ;
      POLYGON 15.800 21.300  15.800 22.300  16.800 22.300  16.800 21.300  
      15.800 21.300  ;
      POLYGON 10.800 3.200  10.800 4.200  11.800 4.200  11.800 3.200  10.800 
      3.200  ;
      POLYGON 10.800 25.300  10.800 26.300  11.800 26.300  11.800 25.300  
      10.800 25.300  ;
      POLYGON 10.800 23.300  10.800 24.300  11.800 24.300  11.800 23.300  
      10.800 23.300  ;
      POLYGON 10.800 21.300  10.800 22.300  11.800 22.300  11.800 21.300  
      10.800 21.300  ;
      POLYGON 7.300 3.200  7.300 4.200  8.300 4.200  8.300 3.200  7.300 3.200  ;
      
      POLYGON 7.300 21.300  7.300 22.300  8.300 22.300  8.300 21.300  7.300 
      21.300  ;
      POLYGON 7.300 23.300  7.300 24.300  8.300 24.300  8.300 23.300  7.300 
      23.300  ;
      POLYGON 7.300 25.300  7.300 26.300  8.300 26.300  8.300 25.300  7.300 
      25.300  ;
      POLYGON 4.300 3.200  4.300 4.200  5.300 4.200  5.300 3.200  4.300 3.200  ;
      
      POLYGON 4.300 25.300  4.300 26.300  5.300 26.300  5.300 25.300  4.300 
      25.300  ;
      POLYGON 4.300 21.300  4.300 22.300  5.300 22.300  5.300 21.300  4.300 
      21.300  ;
      POLYGON 4.300 23.300  4.300 24.300  5.300 24.300  5.300 23.300  4.300 
      23.300  ;
      POLYGON 1.300 25.300  1.300 26.300  2.300 26.300  2.300 25.300  1.300 
      25.300  ;
      POLYGON 1.300 3.200  1.300 4.200  2.300 4.200  2.300 3.200  1.300 3.200  ;
      
      POLYGON 1.300 21.300  1.300 22.300  2.300 22.300  2.300 21.300  1.300 
      21.300  ;
      POLYGON 1.300 23.300  1.300 24.300  2.300 24.300  2.300 23.300  1.300 
      23.300  ;
      POLYGON 27.300 21.300  27.300 22.300  28.300 22.300  28.300 21.300  
      27.300 21.300  ;
      POLYGON 23.800 22.300  23.800 21.300  24.800 21.300  24.800 22.300  
      23.800 22.300  ;
    LAYER FRAME ;
      RECT -0.500 28.500  52.500 30.500  ;
      RECT -0.500 -0.500  52.500 1.500  ;
      POLYGON 0.000 0.000  52.000 0.000  52.000 30.000  0.000 30.000  0.000 
      0.000  ;
    LAYER ML1 ;
      POLYGON 49.300 2.700  51.300 2.700  51.300 4.700  49.300 4.700  49.300 
      2.700  ;
      WIDTH 1.400  ;
      PATH 50.300 22.600 50.300 25.800  ;
      POLYGON 3.300 9.000  3.300 11.000  5.300 11.000  5.300 9.000  3.300 
      9.000  ;
      POLYGON 11.000 9.000  11.000 11.000  13.000 11.000  13.000 9.000  11.000 
      9.000  ;
      POLYGON 21.300 17.700  21.300 19.700  23.300 19.700  23.300 17.700  
      21.300 17.700  ;
      RECT 9.200 -0.500  11.200 1.500  ;
      RECT 26.700 -0.500  28.700 1.500  ;
      RECT 45.000 -0.500  47.000 1.500  ;
      RECT 37.800 5.700  39.800 7.700  ;
      RECT 35.800 13.000  37.800 15.000  ;
      RECT 24.300 17.700  26.300 19.700  ;
      RECT 23.800 5.700  25.800 7.700  ;
      RECT 21.300 9.000  23.300 11.000  ;
      RECT 11.000 9.000  13.000 11.000  ;
      RECT 3.300 9.000  5.300 11.000  ;
      RECT 9.200 28.500  11.200 30.500  ;
      RECT 26.700 28.500  28.700 30.500  ;
      RECT 45.000 28.500  47.000 30.500  ;
      RECT 49.300 24.800  51.300 26.800  ;
      RECT 49.300 22.800  51.300 24.800  ;
      RECT 49.300 20.800  51.300 22.800  ;
      RECT 49.300 2.700  51.300 4.700  ;
      RECT 46.300 24.800  48.300 26.800  ;
      RECT 46.300 22.800  48.300 24.800  ;
      RECT 46.300 20.800  48.300 22.800  ;
      RECT 46.300 2.700  48.300 4.700  ;
      RECT 43.300 24.800  45.300 26.800  ;
      RECT 43.300 22.800  45.300 24.800  ;
      RECT 43.300 20.800  45.300 22.800  ;
      RECT 43.300 2.700  45.300 4.700  ;
      RECT 39.800 2.700  41.800 4.700  ;
      RECT 39.800 24.800  41.800 26.800  ;
      RECT 39.800 22.800  41.800 24.800  ;
      RECT 39.800 20.800  41.800 22.800  ;
      RECT 36.800 2.700  38.800 4.700  ;
      RECT 36.800 24.800  38.800 26.800  ;
      RECT 36.800 22.800  38.800 24.800  ;
      RECT 36.800 20.800  38.800 22.800  ;
      RECT 31.800 2.700  33.800 4.700  ;
      RECT 31.800 24.800  33.800 26.800  ;
      RECT 31.800 22.800  33.800 24.800  ;
      RECT 31.800 20.800  33.800 22.800  ;
      RECT 26.800 2.700  28.800 4.700  ;
      RECT 26.800 22.800  28.800 24.800  ;
      RECT 26.800 24.800  28.800 26.800  ;
      RECT 23.300 2.700  25.300 4.700  ;
      RECT 23.300 24.800  25.300 26.800  ;
      RECT 23.300 22.800  25.300 24.800  ;
      RECT 23.300 20.800  25.300 22.800  ;
      RECT 20.300 2.700  22.300 4.700  ;
      RECT 20.300 24.800  22.300 26.800  ;
      RECT 20.300 22.800  22.300 24.800  ;
      RECT 20.300 20.800  22.300 22.800  ;
      RECT 15.300 2.700  17.300 4.700  ;
      RECT 15.300 22.800  17.300 24.800  ;
      RECT 15.300 24.800  17.300 26.800  ;
      RECT 15.300 20.800  17.300 22.800  ;
      RECT 10.300 2.700  12.300 4.700  ;
      RECT 10.300 24.800  12.300 26.800  ;
      RECT 10.300 22.800  12.300 24.800  ;
      RECT 10.300 20.800  12.300 22.800  ;
      RECT 6.800 2.700  8.800 4.700  ;
      RECT 6.800 20.800  8.800 22.800  ;
      RECT 6.800 22.800  8.800 24.800  ;
      RECT 6.800 24.800  8.800 26.800  ;
      RECT 3.800 2.700  5.800 4.700  ;
      RECT 3.800 24.800  5.800 26.800  ;
      RECT 3.800 20.800  5.800 22.800  ;
      RECT 3.800 22.800  5.800 24.800  ;
      RECT 0.800 24.800  2.800 26.800  ;
      RECT 0.800 2.700  2.800 4.700  ;
      RECT 0.800 20.800  2.800 22.800  ;
      RECT 0.800 22.800  2.800 24.800  ;
      POLYGON -0.500 30.500  -0.500 28.500  4.100 28.500  4.100 21.900  5.500 
      21.900  5.500 28.500  10.600 28.500  10.600 21.900  12.000 21.900  
      12.000 28.500  20.600 28.500  20.600 21.900  22.000 21.900  22.000 
      28.500  27.100 28.500  27.100 21.100  28.500 21.100  28.500 28.500  
      37.100 28.500  37.100 21.900  38.500 21.900  38.500 28.500  46.600 
      28.500  46.600 21.900  48.000 21.900  48.000 28.500  52.500 28.500  
      52.500 30.500  -0.500 30.500  ;
      RECT 26.800 20.800  28.800 22.800  ;
      POLYGON -0.500 1.500  -0.500 -0.500  52.500 -0.500  52.500 1.500  48.000 
      1.500  48.000 4.400  46.600 4.400  46.600 1.500  38.500 1.500  38.500 
      4.400  37.100 4.400  37.100 1.500  28.500 1.500  28.500 4.400  27.100 
      4.400  27.100 1.500  22.000 1.500  22.000 4.400  20.600 4.400  20.600 
      1.500  12.000 1.500  12.000 4.400  10.600 4.400  10.600 1.500  5.500 
      1.500  5.500 4.400  4.100 4.400  4.100 1.500  -0.500 1.500  ;
      POLYGON 1.100 26.500  1.100 21.900  1.300 21.900  1.300 3.000  2.300 
      3.000  2.300 6.200  4.800 6.200  4.800 5.700  6.800 5.700  6.800 7.700  
      4.800 7.700  4.800 7.200  2.300 7.200  2.300 12.500  4.300 12.500  4.300 
      12.000  6.300 12.000  6.300 14.000  4.300 14.000  4.300 13.500  2.300 
      13.500  2.300 18.300  4.800 18.300  4.800 17.800  6.800 17.800  6.800 
      19.800  4.800 19.800  4.800 19.300  2.300 19.300  2.300 21.900  2.500 
      21.900  2.500 26.500  1.100 26.500  ;
      POLYGON 7.300 16.700  7.300 9.000  7.800 9.000  7.800 3.000  8.800 3.000 
       8.800 6.200  13.800 6.200  13.800 5.700  15.800 5.700  15.800 7.700  
      13.800 7.700  13.800 7.200  8.800 7.200  8.800 10.000  8.300 10.000  
      8.300 15.700  16.300 15.700  16.300 15.000  18.300 15.000  18.300 15.700 
       32.800 15.700  32.800 17.700  30.800 17.700  30.800 16.700  18.300 
      16.700  18.300 17.000  16.300 17.000  16.300 16.700  8.800 16.700  8.800 
      26.500  7.800 26.500  7.800 16.700  7.300 16.700  ;
      POLYGON 15.800 4.700  15.800 3.200  16.800 3.200  16.800 3.700  17.300 
      3.700  17.300 9.500  21.300 9.500  21.300 9.000  23.300 9.000  23.300 
      11.000  21.300 11.000  21.300 10.500  16.300 10.500  16.300 4.700  
      15.800 4.700  ;
      POLYGON 15.600 26.500  15.600 21.900  15.800 21.900  15.800 18.300  
      21.300 18.300  21.300 17.700  23.300 17.700  23.300 19.700  21.300 
      19.700  21.300 19.300  16.800 19.300  16.800 21.900  17.000 21.900  
      17.000 26.500  15.600 26.500  ;
      POLYGON 9.300 14.000  9.300 12.000  11.300 12.000  11.300 12.500  14.300 
      12.500  14.300 12.000  16.300 12.000  16.300 12.500  27.800 12.500  
      27.800 12.000  29.800 12.000  29.800 12.500  34.500 12.500  34.500 
      12.700  34.800 12.700  34.800 14.700  32.800 14.700  32.800 13.500  
      29.800 13.500  29.800 14.000  27.800 14.000  27.800 13.500  16.300 
      13.500  16.300 14.000  14.300 14.000  14.300 13.500  11.300 13.500  
      11.300 14.000  9.300 14.000  ;
      POLYGON 19.300 7.700  19.300 5.700  21.300 5.700  21.300 6.200  23.800 
      6.200  23.800 2.900  24.800 2.900  24.800 5.700  25.800 5.700  25.800 
      7.700  23.800 7.700  23.800 7.200  21.300 7.200  21.300 7.700  19.300 
      7.700  ;
      POLYGON 24.300 19.700  24.300 17.700  26.300 17.700  26.300 19.700  
      25.500 19.700  25.500 22.300  25.000 22.300  25.000 26.500  23.600 
      26.500  23.600 21.100  24.500 21.100  24.500 19.700  24.300 19.700  ;
      POLYGON 32.100 26.500  32.100 21.900  32.300 21.900  32.300 18.700  
      37.800 18.700  37.800 17.700  39.800 17.700  39.800 19.700  33.300 
      19.700  33.300 21.900  33.500 21.900  33.500 26.500  32.100 26.500  ;
      POLYGON 37.800 19.700  37.800 17.700  39.800 17.700  39.800 19.700  
      37.800 19.700  ;
      POLYGON 36.300 14.500  36.300 13.500  40.800 13.500  40.800 3.200  
      41.800 3.200  41.800 8.200  44.300 8.200  44.300 7.700  46.300 7.700  
      46.300 9.700  44.300 9.700  44.300 9.200  41.800 9.200  41.800 16.700  
      44.300 16.700  44.300 16.200  46.300 16.200  46.300 18.200  44.300 
      18.200  44.300 17.700  41.800 17.700  41.800 26.300  40.800 26.300  
      40.800 14.500  36.300 14.500  ;
      POLYGON 43.800 6.700  43.800 3.000  44.800 3.000  44.800 5.700  49.300 
      5.700  49.300 7.700  48.500 7.700  48.500 17.900  49.300 17.900  49.300 
      19.900  44.700 19.900  44.700 21.900  45.000 21.900  45.000 26.500  
      43.600 26.500  43.600 21.900  43.700 21.900  43.700 18.900  47.300 
      18.900  47.300 17.900  47.500 17.900  47.500 7.700  47.300 7.700  47.300 
      6.700  43.800 6.700  ;
      POLYGON 49.500 12.500  49.500 10.500  50.300 10.500  50.300 2.700  
      51.300 2.700  51.300 10.500  51.500 10.500  51.500 12.500  51.300 12.500 
       51.300 26.500  50.300 26.500  50.300 12.500  49.500 12.500  ;
      POLYGON 32.300 7.200  32.300 3.200  33.300 3.200  33.300 6.200  37.800 
      6.200  37.800 5.700  39.800 5.700  39.800 7.700  37.800 7.700  37.800 
      7.200  32.300 7.200  ;
    LAYER ML2 ;
      POLYGON 11.000 9.000  11.000 11.000  13.000 11.000  13.000 9.000  11.000 
      9.000  ;
      POLYGON 3.300 11.000  3.300 9.000  5.300 9.000  5.300 11.000  3.300 
      11.000  ;
      POLYGON 21.300 11.000  21.300 9.000  23.300 9.000  23.300 11.000  22.800 
      11.000  22.800 17.700  23.300 17.700  23.300 19.700  21.300 19.700  
      21.300 17.700  21.800 17.700  21.800 11.000  21.300 11.000  ;
      POLYGON 23.800 7.700  23.800 5.700  25.800 5.700  25.800 7.700  25.300 
      7.700  25.300 17.700  26.300 17.700  26.300 19.700  24.300 19.700  
      24.300 7.700  23.800 7.700  ;
      POLYGON 37.800 7.700  37.800 5.700  39.800 5.700  39.800 7.700  39.300 
      7.700  39.300 17.700  39.800 17.700  39.800 19.700  37.800 19.700  
      37.800 17.700  38.300 17.700  38.300 7.700  37.800 7.700  ;
      POLYGON 49.500 12.500  49.500 10.500  51.500 10.500  51.500 12.500  
      49.500 12.500  ;
    LAYER POL ;
      WIDTH 1.000  ;
      PATH 6.300 18.600 6.300 27.300  ;
      POLYGON 4.800 17.800  4.800 19.800  6.800 19.800  6.800 17.800  4.800 
      17.800  ;
      POLYGON 4.800 7.700  4.800 5.700  5.800 5.700  5.800 1.700  6.800 1.700  
      6.800 7.700  4.800 7.700  ;
      POLYGON 2.800 27.800  2.800 1.700  3.800 1.700  3.800 9.000  5.300 9.000 
       5.300 11.000  3.800 11.000  3.800 27.800  2.800 27.800  ;
      POLYGON 4.300 14.000  4.300 12.000  6.300 12.000  6.300 12.500  9.300 
      12.500  9.300 12.000  11.300 12.000  11.300 14.000  9.300 14.000  9.300 
      13.500  6.300 13.500  6.300 14.000  4.300 14.000  ;
      POLYGON 11.000 11.000  11.000 9.000  12.300 9.000  12.300 1.900  13.300 
      1.900  13.300 27.600  12.300 27.600  12.300 11.000  11.000 11.000  ;
      POLYGON 13.800 7.700  13.800 5.700  14.300 5.700  14.300 1.900  15.300 
      1.900  15.300 5.700  15.800 5.700  15.800 7.700  13.800 7.700  ;
      POLYGON 21.300 19.700  21.300 17.700  23.300 17.700  23.300 27.600  
      22.300 27.600  22.300 19.700  21.300 19.700  ;
      POLYGON 16.300 17.000  16.300 15.000  18.300 15.000  18.300 27.600  
      17.300 27.600  17.300 17.000  16.300 17.000  ;
      POLYGON 14.300 27.600  14.300 12.000  15.300 12.000  15.300 11.000  
      17.300 11.000  17.300 1.900  18.300 1.900  18.300 12.000  16.300 12.000  
      16.300 14.000  15.300 14.000  15.300 27.600  14.300 27.600  ;
      POLYGON 19.300 27.500  19.300 1.800  20.300 1.800  20.300 5.700  21.300 
      5.700  21.300 7.700  20.300 7.700  20.300 27.500  19.300 27.500  ;
      POLYGON 21.300 11.000  21.300 9.000  22.300 9.000  22.300 1.900  23.300 
      1.900  23.300 11.000  21.300 11.000  ;
      POLYGON 23.800 7.700  23.800 5.700  24.800 5.700  24.800 5.200  28.800 
      5.200  28.800 1.900  29.800 1.900  29.800 6.200  25.800 6.200  25.800 
      7.700  23.800 7.700  ;
      POLYGON 24.300 19.700  24.300 17.700  26.300 17.700  26.300 18.700  
      29.800 18.700  29.800 27.600  28.800 27.600  28.800 19.700  24.300 
      19.700  ;
      POLYGON 27.800 14.000  27.800 12.000  28.300 12.000  28.300 7.200  
      30.800 7.200  30.800 1.900  31.800 1.900  31.800 8.200  29.300 8.200  
      29.300 12.000  29.800 12.000  29.800 14.000  27.800 14.000  ;
      POLYGON 30.800 27.600  30.800 10.700  33.800 10.700  33.800 1.900  
      34.800 1.900  34.800 11.700  31.800 11.700  31.800 15.700  32.800 15.700 
       32.800 17.700  31.800 17.700  31.800 27.600  30.800 27.600  ;
      POLYGON 37.800 7.700  37.800 5.700  38.800 5.700  38.800 1.900  39.800 
      1.900  39.800 7.700  37.800 7.700  ;
      POLYGON 35.800 27.600  35.800 1.900  36.800 1.900  36.800 13.000  37.800 
      13.000  37.800 15.000  36.800 15.000  36.800 27.600  35.800 27.600  ;
      POLYGON 32.800 14.700  32.800 12.700  34.800 12.700  34.800 27.600  
      33.800 27.600  33.800 14.700  32.800 14.700  ;
      POLYGON 37.800 19.700  37.800 17.700  39.800 17.700  39.800 27.600  
      38.800 27.600  38.800 19.700  37.800 19.700  ;
      POLYGON 44.300 18.200  44.300 16.200  46.300 16.200  46.300 27.600  
      45.300 27.600  45.300 18.200  44.300 18.200  ;
      POLYGON 47.300 19.900  47.300 17.900  49.300 17.900  49.300 27.600  
      48.300 27.600  48.300 19.900  47.300 19.900  ;
      POLYGON 47.300 7.700  47.300 5.700  48.300 5.700  48.300 1.900  49.300 
      1.900  49.300 7.700  47.300 7.700  ;
      POLYGON 44.300 9.700  44.300 7.700  45.300 7.700  45.300 1.900  46.300 
      1.900  46.300 9.700  44.300 9.700  ;
    LAYER VIA1 ;
      POLYGON 38.300 18.200  38.300 19.200  39.300 19.200  39.300 18.200  
      38.300 18.200  ;
      POLYGON 38.300 6.200  38.300 7.200  39.300 7.200  39.300 6.200  38.300 
      6.200  ;
      POLYGON 24.800 18.200  24.800 19.200  25.800 19.200  25.800 18.200  
      24.800 18.200  ;
      POLYGON 24.300 6.200  24.300 7.200  25.300 7.200  25.300 6.200  24.300 
      6.200  ;
      POLYGON 21.800 9.500  21.800 10.500  22.800 10.500  22.800 9.500  21.800 
      9.500  ;
      POLYGON 21.800 18.200  21.800 19.200  22.800 19.200  22.800 18.200  
      21.800 18.200  ;
      POLYGON 11.500 9.500  11.500 10.500  12.500 10.500  12.500 9.500  11.500 
      9.500  ;
      POLYGON 3.800 9.500  3.800 10.500  4.800 10.500  4.800 9.500  3.800 
      9.500  ;
      POLYGON 50.000 11.000  50.000 12.000  51.000 12.000  51.000 11.000  
      50.000 11.000  ;
  END
END dff1m2LEF


END LIBRARY
