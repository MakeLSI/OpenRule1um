VERSION 5.3 ;

NAMESCASESENSITIVE ON ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS











MACRO cinvLEF
  CLASS BLOCK ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER POL ;
        POLYGON 6.500 13.500  6.500 11.500  7.800 11.500  7.800 1.700  8.800 
        1.700  8.800 26.500  7.800 26.500  7.800 13.500  6.500 13.500  ;
    END
    PORT
      LAYER ML1 ;
        POLYGON 6.500 11.500  6.500 13.500  8.500 13.500  8.500 11.500  6.500 
        11.500  ;
    END
  END A
  PIN OE
    DIRECTION INPUT ;
    PORT
      LAYER POL ;
        POLYGON 1.000 16.500  1.000 14.500  2.000 14.500  2.000 6.000  2.800 
        6.000  2.800 1.700  3.800 1.700  3.800 6.000  5.800 6.000  5.800 1.700 
         6.800 1.700  6.800 7.000  3.000 7.000  3.000 15.000  3.800 15.000  
        3.800 26.500  2.800 26.500  2.800 16.500  1.000 16.500  ;
    END
    PORT
      LAYER ML1 ;
        POLYGON 1.000 14.500  1.000 16.500  3.000 16.500  3.000 14.500  1.000 
        14.500  ;
    END
  END OE
  PIN VDD
    DIRECTION INOUT ;
    PORT
      LAYER ML1 ;
        POLYGON -0.500 30.500  -0.500 28.500  4.100 28.500  4.100 20.600  
        5.500 20.600  5.500 28.500  12.000 28.500  12.000 30.500  -0.500 
        30.500  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    PORT
      LAYER ML1 ;
        POLYGON -0.500 1.500  -0.500 -0.500  12.000 -0.500  12.000 1.500  
        5.300 1.500  5.300 4.200  4.300 4.200  4.300 1.500  -0.500 1.500  ;
    END
  END VSS
  PIN YB
    DIRECTION OUTPUT ;
    PORT
      LAYER ML1 ;
        POLYGON 9.000 9.200  9.000 7.200  9.300 7.200  9.300 3.200  10.300 
        3.200  10.300 7.200  11.000 7.200  11.000 9.200  10.500 9.200  10.500 
        18.500  10.300 18.500  10.300 20.600  10.500 20.600  10.500 25.200  
        9.100 25.200  9.100 20.600  9.300 20.600  9.300 17.500  9.500 17.500  
        9.500 9.200  9.000 9.200  ;
    END
  END YB
  OBS
    LAYER CNT ;
      POLYGON 4.300 24.000  4.300 25.000  5.300 25.000  5.300 24.000  4.300 
      24.000  ;
      POLYGON 4.300 3.200  4.300 4.200  5.300 4.200  5.300 3.200  4.300 3.200  ;
      
      POLYGON 9.300 3.200  9.300 4.200  10.300 4.200  10.300 3.200  9.300 
      3.200  ;
      POLYGON 9.300 20.000  9.300 21.000  10.300 21.000  10.300 20.000  9.300 
      20.000  ;
      POLYGON 9.300 22.000  9.300 23.000  10.300 23.000  10.300 22.000  9.300 
      22.000  ;
      POLYGON 9.300 24.000  9.300 25.000  10.300 25.000  10.300 24.000  9.300 
      24.000  ;
      POLYGON 5.300 15.000  5.300 16.000  6.300 16.000  6.300 15.000  5.300 
      15.000  ;
      POLYGON 7.000 12.000  7.000 13.000  8.000 13.000  8.000 12.000  7.000 
      12.000  ;
      POLYGON 6.500 29.000  6.500 30.000  7.500 30.000  7.500 29.000  6.500 
      29.000  ;
      POLYGON 1.500 15.000  1.500 16.000  2.500 16.000  2.500 15.000  1.500 
      15.000  ;
      POLYGON 5.500 0.000  5.500 1.000  6.500 1.000  6.500 0.000  5.500 0.000  ;
      
      POLYGON 4.300 20.000  4.300 21.000  5.300 21.000  5.300 20.000  4.300 
      20.000  ;
      POLYGON 4.300 22.000  4.300 23.000  5.300 23.000  5.300 22.000  4.300 
      22.000  ;
      POLYGON 1.300 24.000  1.300 25.000  2.300 25.000  2.300 24.000  1.300 
      24.000  ;
      POLYGON 1.300 3.200  1.300 4.200  2.300 4.200  2.300 3.200  1.300 3.200  ;
      
      POLYGON 1.300 20.000  1.300 21.000  2.300 21.000  2.300 20.000  1.300 
      20.000  ;
      POLYGON 1.300 22.000  1.300 23.000  2.300 23.000  2.300 22.000  1.300 
      22.000  ;
    LAYER FRAME ;
      RECT -0.500 28.500  12.000 30.500  ;
      RECT -0.500 -0.500  12.000 1.500  ;
      POLYGON 0.000 0.000  11.500 0.000  11.500 30.000  0.000 30.000  0.000 
      0.000  ;
    LAYER ML1 ;
      RECT 5.000 -0.500  7.000 1.500  ;
      POLYGON 1.000 14.500  1.000 16.500  3.000 16.500  3.000 14.500  1.000 
      14.500  ;
      WIDTH 1.400  ;
      PATH 1.800 21.300 1.800 24.500  ;
      POLYGON 6.500 11.500  6.500 13.500  8.500 13.500  8.500 11.500  6.500 
      11.500  ;
      RECT 1.000 14.500  3.000 16.500  ;
      RECT 6.000 28.500  8.000 30.500  ;
      RECT 6.500 11.500  8.500 13.500  ;
      RECT 8.800 23.500  10.800 25.500  ;
      RECT 8.800 21.500  10.800 23.500  ;
      RECT 8.800 19.500  10.800 21.500  ;
      RECT 8.800 2.700  10.800 4.700  ;
      RECT 3.800 2.700  5.800 4.700  ;
      RECT 3.800 23.500  5.800 25.500  ;
      RECT 3.800 19.500  5.800 21.500  ;
      RECT 3.800 21.500  5.800 23.500  ;
      RECT 0.800 23.500  2.800 25.500  ;
      RECT 0.800 2.700  2.800 4.700  ;
      RECT 0.800 19.500  2.800 21.500  ;
      RECT 0.800 21.500  2.800 23.500  ;
      POLYGON -0.500 30.500  -0.500 28.500  4.100 28.500  4.100 20.600  5.500 
      20.600  5.500 28.500  12.000 28.500  12.000 30.500  -0.500 30.500  ;
      POLYGON -0.500 1.500  -0.500 -0.500  12.000 -0.500  12.000 1.500  5.300 
      1.500  5.300 4.200  4.300 4.200  4.300 1.500  -0.500 1.500  ;
      POLYGON 1.300 8.500  1.300 3.200  2.300 3.200  2.300 7.500  5.500 7.500  
      5.500 14.500  6.800 14.500  6.800 16.500  5.500 16.500  5.500 18.500  
      2.300 18.500  2.300 25.000  1.300 25.000  1.300 17.500  4.500 17.500  
      4.500 8.500  1.300 8.500  ;
      POLYGON 9.000 9.200  9.000 7.200  9.300 7.200  9.300 3.200  10.300 3.200 
       10.300 7.200  11.000 7.200  11.000 9.200  10.500 9.200  10.500 18.500  
      10.300 18.500  10.300 20.600  10.500 20.600  10.500 25.200  9.100 25.200 
       9.100 20.600  9.300 20.600  9.300 17.500  9.500 17.500  9.500 9.200  
      9.000 9.200  ;
    LAYER ML2 ;
      POLYGON 9.000 9.200  9.000 7.200  11.000 7.200  11.000 9.200  9.000 
      9.200  ;
      POLYGON 6.500 11.500  6.500 13.500  8.500 13.500  8.500 11.500  6.500 
      11.500  ;
      POLYGON 1.000 14.500  1.000 16.500  3.000 16.500  3.000 14.500  1.000 
      14.500  ;
    LAYER POL ;
      POLYGON 6.500 13.500  6.500 11.500  7.800 11.500  7.800 1.700  8.800 
      1.700  8.800 26.500  7.800 26.500  7.800 13.500  6.500 13.500  ;
      POLYGON 4.800 16.500  4.800 14.500  6.800 14.500  6.800 26.500  5.800 
      26.500  5.800 16.500  4.800 16.500  ;
      POLYGON 1.000 16.500  1.000 14.500  2.000 14.500  2.000 6.000  2.800 
      6.000  2.800 1.700  3.800 1.700  3.800 6.000  5.800 6.000  5.800 1.700  
      6.800 1.700  6.800 7.000  3.000 7.000  3.000 15.000  3.800 15.000  3.800 
      26.500  2.800 26.500  2.800 16.500  1.000 16.500  ;
    LAYER VIA1 ;
      POLYGON 7.000 12.000  7.000 13.000  8.000 13.000  8.000 12.000  7.000 
      12.000  ;
      POLYGON 9.500 7.700  9.500 8.700  10.500 8.700  10.500 7.700  9.500 
      7.700  ;
      POLYGON 1.500 15.000  1.500 16.000  2.500 16.000  2.500 15.000  1.500 
      15.000  ;
  END
END cinvLEF


END LIBRARY
