VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO or31
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 15.500 BY 30.000 ;
  SYMMETRY X Y ;
  SITE unit ;
 
  PIN A
    USE SIGNAL ;
    PORT
      LAYER ML1 ;
        POLYGON 1.000 14.500  1.000 16.500  3.000 16.500  3.000 14.500  1.000 
        14.500  ;
    END
    PORT
      LAYER ML2 ;
        POLYGON 1.000 14.500  1.000 16.500  3.000 16.500  3.000 14.500  1.000 
        14.500  ;
    END
  END A
  PIN B
    USE SIGNAL ;
    PORT
      LAYER ML2 ;
        POLYGON 4.000 11.500  4.000 13.500  6.000 13.500  6.000 11.500  4.000 
        11.500  ;
    END
    PORT
      LAYER ML1 ;
        POLYGON 4.000 11.500  4.000 13.500  6.000 13.500  6.000 11.500  4.000 
        11.500  ;
    END
  END B
  PIN C
    USE SIGNAL ;
    PORT
      LAYER ML1 ;
        POLYGON 7.000 12.000  7.000 14.000  9.000 14.000  9.000 12.000  7.000 
        12.000  ;
    END
    PORT
      LAYER ML2 ;
        POLYGON 7.000 12.000  7.000 14.000  9.000 14.000  9.000 12.000  7.000 
        12.000  ;
    END
  END C
  PIN VDD
    USE POWER ;
    PORT
      LAYER ML1 ;
        RECT -0.500 28.500  16.000 30.500  ;
    END
  END VDD
  PIN VSS
    USE GROUND ;
    PORT
      LAYER ML1 ;
        RECT -0.500 -0.500  16.000 1.500  ;
    END
  END VSS
  PIN Y
    USE SIGNAL ;
    PORT
      LAYER ML2 ;
        RECT 13.000 9.000  15.000 11.000  ;
    END
    PORT
      LAYER ML1 ;
        RECT 13.000 9.000  15.000 11.000  ;
    END
    PORT
      LAYER ML1 ;
        WIDTH 1.000  ;
        PATH 13.800 3.900 13.800 16.500 12.800 16.500 12.800 20.500  ;
    END
  END Y
  OBS

    LAYER ML1 ;

      WIDTH 1.400  ;
      PATH 2.800 21.300 2.800 24.500  ;
      WIDTH 1.000  ;
      PATH 4.800 1.000 4.800 3.800  ;

      WIDTH 1.000  ;
      PATH 2.800 20.500 2.800 18.000 10.500 18.000 10.500 8.000 1.800 8.000 
      1.800 3.800  ;

      WIDTH 1.000  ;
      PATH 7.800 3.900 7.800 8.000  ;

      WIDTH 1.400  ;
      PATH 9.800 21.300 9.800 28.500  ;
      WIDTH 1.000  ;
      PATH 10.800 1.000 10.800 3.800  ;
      WIDTH 1.400  ;
      PATH 12.800 21.300 12.800 24.500  ;
      WIDTH 1.000  ;
      PATH 13.800 3.900 13.800 16.500 12.800 16.500 12.800 20.500  ;

    VIA 1.800 3.800  dcont ;
    VIA 2.800 24.500  dcont ;
    VIA 2.800 20.500  dcont ;
    VIA 2.800 22.500  dcont ;
    VIA 4.800 3.800  dcont ;
    VIA 7.800 3.800  dcont ;
    VIA 9.800 24.500  dcont ;
    VIA 9.800 22.500  dcont ;
    VIA 9.800 20.500  dcont ;
    VIA 10.800 3.800  dcont ;
    VIA 12.800 24.500  dcont ;
    VIA 12.800 22.500  dcont ;
    VIA 12.800 20.500  dcont ;
    VIA 13.800 3.800  dcont ;
    VIA 5.000 12.500  pcont ;
    VIA 8.200 29.500  nsubcont ;
    VIA 8.000 13.000  pcont ;
    VIA 11.300 13.000  pcont ;
    VIA 2.000 15.500  pcont ;
    VIA 6.500 0.500  psubcont ;
  END
END or31

MACRO dcont
  CLASS CORE ;
  OBS
    LAYER ML1 ;
      RECT -1.000 -1.000  1.000 1.000  ;
  END
END dcont

MACRO pcont
  CLASS CORE ;
  OBS
    LAYER ML1 ;
      RECT -1.000 -1.000  1.000 1.000  ;
  END
END pcont

MACRO nsubcont
  CLASS CORE ;
  OBS
    LAYER ML1 ;
      RECT -1.000 -1.000  1.000 1.000  ;
  END
END nsubcont

MACRO psubcont
  CLASS CORE ;
  OBS
    LAYER ML1 ;
      RECT -1.000 -1.000  1.000 1.000  ;
  END
END psubcont


END LIBRARY
