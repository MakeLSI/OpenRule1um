VERSION 5.3 ;

NAMESCASESENSITIVE ON ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS











MACRO sff1m2LEF
  CLASS BLOCK ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER POL ;
        POLYGON 2.800 27.800  2.800 1.700  3.800 1.700  3.800 9.000  5.500 
        9.000  5.500 11.000  3.800 11.000  3.800 27.800  2.800 27.800  ;
    END
    PORT
      LAYER ML1 ;
        POLYGON 3.500 9.000  3.500 11.000  5.500 11.000  5.500 9.000  3.500 
        9.000  ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER POL ;
        POLYGON 11.000 11.000  11.000 9.000  12.300 9.000  12.300 1.900  
        13.300 1.900  13.300 27.600  12.300 27.600  12.300 11.000  11.000 
        11.000  ;
    END
    PORT
      LAYER ML1 ;
        POLYGON 11.000 9.000  11.000 11.000  13.000 11.000  13.000 9.000  
        11.000 9.000  ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER ML1 ;
        POLYGON 53.500 12.500  53.500 10.500  54.300 10.500  54.300 2.700  
        55.300 2.700  55.300 10.500  55.500 10.500  55.500 12.500  55.300 
        12.500  55.300 26.500  54.300 26.500  54.300 12.500  53.500 12.500  ;
    END
  END Q
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER POL ;
        POLYGON 41.300 27.600  41.300 11.500  42.800 11.500  42.800 1.900  
        43.800 1.900  43.800 10.500  45.000 10.500  45.000 12.500  42.300 
        12.500  42.300 27.600  41.300 27.600  ;
    END
    PORT
      LAYER ML1 ;
        POLYGON 43.000 10.500  43.000 12.500  45.000 12.500  45.000 10.500  
        43.000 10.500  ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    PORT
      LAYER ML1 ;
        POLYGON -0.500 30.500  -0.500 28.500  4.100 28.500  4.100 21.900  
        5.500 21.900  5.500 28.500  10.600 28.500  10.600 21.900  12.000 
        21.900  12.000 28.500  20.600 28.500  20.600 21.900  22.000 21.900  
        22.000 28.500  26.600 28.500  26.600 23.100  28.000 23.100  28.000 
        28.500  36.600 28.500  36.600 21.900  38.000 21.900  38.000 28.500  
        42.600 28.500  42.600 21.900  44.000 21.900  44.000 28.500  50.600 
        28.500  50.600 21.900  52.000 21.900  52.000 28.500  56.500 28.500  
        56.500 30.500  -0.500 30.500  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    PORT
      LAYER ML1 ;
        POLYGON -0.500 1.500  -0.500 -0.500  56.500 -0.500  56.500 1.500  
        52.000 1.500  52.000 4.400  50.600 4.400  50.600 1.500  40.500 1.500  
        40.500 4.400  39.100 4.400  39.100 1.500  30.500 1.500  30.500 4.400  
        29.100 4.400  29.100 1.500  22.000 1.500  22.000 4.400  20.600 4.400  
        20.600 1.500  12.000 1.500  12.000 4.400  10.600 4.400  10.600 1.500  
        5.500 1.500  5.500 4.400  4.100 4.400  4.100 1.500  -0.500 1.500  ;
    END
  END VSS
  OBS
    LAYER CNT ;
      POLYGON 37.800 13.500  37.800 14.500  38.800 14.500  38.800 13.500  
      37.800 13.500  ;
      POLYGON 37.800 18.200  37.800 19.200  38.800 19.200  38.800 18.200  
      37.800 18.200  ;
      POLYGON 40.300 6.200  40.300 7.200  41.300 7.200  41.300 6.200  40.300 
      6.200  ;
      POLYGON 43.500 11.000  43.500 12.000  44.500 12.000  44.500 11.000  
      43.500 11.000  ;
      POLYGON 48.800 8.200  48.800 9.200  49.800 9.200  49.800 8.200  48.800 
      8.200  ;
      POLYGON 48.800 16.700  48.800 17.700  49.800 17.700  49.800 16.700  
      48.800 16.700  ;
      POLYGON 51.800 6.200  51.800 7.200  52.800 7.200  52.800 6.200  51.800 
      6.200  ;
      POLYGON 51.800 18.400  51.800 19.400  52.800 19.400  52.800 18.400  
      51.800 18.400  ;
      POLYGON 49.500 0.000  49.500 1.000  50.500 1.000  50.500 0.000  49.500 
      0.000  ;
      POLYGON 27.200 0.000  27.200 1.000  28.200 1.000  28.200 0.000  27.200 
      0.000  ;
      POLYGON 9.700 0.000  9.700 1.000  10.700 1.000  10.700 0.000  9.700 
      0.000  ;
      POLYGON 32.800 13.200  32.800 14.200  33.800 14.200  33.800 13.200  
      32.800 13.200  ;
      POLYGON 30.800 16.200  30.800 17.200  31.800 17.200  31.800 16.200  
      30.800 16.200  ;
      POLYGON 27.800 12.500  27.800 13.500  28.800 13.500  28.800 12.500  
      27.800 12.500  ;
      POLYGON 27.800 18.200  27.800 19.200  28.800 19.200  28.800 18.200  
      27.800 18.200  ;
      POLYGON 26.800 6.200  26.800 7.200  27.800 7.200  27.800 6.200  26.800 
      6.200  ;
      POLYGON 24.800 9.500  24.800 10.500  25.800 10.500  25.800 9.500  24.800 
      9.500  ;
      POLYGON 21.800 9.500  21.800 10.500  22.800 10.500  22.800 9.500  21.800 
      9.500  ;
      POLYGON 21.800 18.200  21.800 19.200  22.800 19.200  22.800 18.200  
      21.800 18.200  ;
      POLYGON 19.800 6.200  19.800 7.200  20.800 7.200  20.800 6.200  19.800 
      6.200  ;
      POLYGON 16.800 15.500  16.800 16.500  17.800 16.500  17.800 15.500  
      16.800 15.500  ;
      POLYGON 14.800 12.500  14.800 13.500  15.800 13.500  15.800 12.500  
      14.800 12.500  ;
      POLYGON 14.300 6.200  14.300 7.200  15.300 7.200  15.300 6.200  14.300 
      6.200  ;
      POLYGON 11.500 9.500  11.500 10.500  12.500 10.500  12.500 9.500  11.500 
      9.500  ;
      POLYGON 9.800 12.500  9.800 13.500  10.800 13.500  10.800 12.500  9.800 
      12.500  ;
      POLYGON 5.300 6.200  5.300 7.200  6.300 7.200  6.300 6.200  5.300 6.200  ;
      
      POLYGON 5.300 18.300  5.300 19.300  6.300 19.300  6.300 18.300  5.300 
      18.300  ;
      POLYGON 4.800 12.500  4.800 13.500  5.800 13.500  5.800 12.500  4.800 
      12.500  ;
      POLYGON 4.000 9.500  4.000 10.500  5.000 10.500  5.000 9.500  4.000 
      9.500  ;
      POLYGON 9.700 29.000  9.700 30.000  10.700 30.000  10.700 29.000  9.700 
      29.000  ;
      POLYGON 27.200 29.000  27.200 30.000  28.200 30.000  28.200 29.000  
      27.200 29.000  ;
      POLYGON 49.500 29.000  49.500 30.000  50.500 30.000  50.500 29.000  
      49.500 29.000  ;
      POLYGON 53.800 25.300  53.800 26.300  54.800 26.300  54.800 25.300  
      53.800 25.300  ;
      POLYGON 53.800 23.300  53.800 24.300  54.800 24.300  54.800 23.300  
      53.800 23.300  ;
      POLYGON 53.800 21.300  53.800 22.300  54.800 22.300  54.800 21.300  
      53.800 21.300  ;
      POLYGON 53.800 3.200  53.800 4.200  54.800 4.200  54.800 3.200  53.800 
      3.200  ;
      POLYGON 50.800 25.300  50.800 26.300  51.800 26.300  51.800 25.300  
      50.800 25.300  ;
      POLYGON 50.800 23.300  50.800 24.300  51.800 24.300  51.800 23.300  
      50.800 23.300  ;
      POLYGON 50.800 21.300  50.800 22.300  51.800 22.300  51.800 21.300  
      50.800 21.300  ;
      POLYGON 50.800 3.200  50.800 4.200  51.800 4.200  51.800 3.200  50.800 
      3.200  ;
      POLYGON 47.800 25.300  47.800 26.300  48.800 26.300  48.800 25.300  
      47.800 25.300  ;
      POLYGON 47.800 23.300  47.800 24.300  48.800 24.300  48.800 23.300  
      47.800 23.300  ;
      POLYGON 47.800 21.300  47.800 22.300  48.800 22.300  48.800 21.300  
      47.800 21.300  ;
      POLYGON 47.800 3.200  47.800 4.200  48.800 4.200  48.800 3.200  47.800 
      3.200  ;
      POLYGON 44.300 3.200  44.300 4.200  45.300 4.200  45.300 3.200  44.300 
      3.200  ;
      POLYGON 42.800 21.300  42.800 22.300  43.800 22.300  43.800 21.300  
      42.800 21.300  ;
      POLYGON 42.800 23.300  42.800 24.300  43.800 24.300  43.800 23.300  
      42.800 23.300  ;
      POLYGON 42.800 25.300  42.800 26.300  43.800 26.300  43.800 25.300  
      42.800 25.300  ;
      POLYGON 39.800 25.300  39.800 26.300  40.800 26.300  40.800 25.300  
      39.800 25.300  ;
      POLYGON 39.800 23.300  39.800 24.300  40.800 24.300  40.800 23.300  
      39.800 23.300  ;
      POLYGON 39.800 21.300  39.800 22.300  40.800 22.300  40.800 21.300  
      39.800 21.300  ;
      POLYGON 39.300 3.200  39.300 4.200  40.300 4.200  40.300 3.200  39.300 
      3.200  ;
      POLYGON 36.800 25.300  36.800 26.300  37.800 26.300  37.800 25.300  
      36.800 25.300  ;
      POLYGON 36.800 23.300  36.800 24.300  37.800 24.300  37.800 23.300  
      36.800 23.300  ;
      POLYGON 36.800 21.300  36.800 22.300  37.800 22.300  37.800 21.300  
      36.800 21.300  ;
      POLYGON 34.300 3.200  34.300 4.200  35.300 4.200  35.300 3.200  34.300 
      3.200  ;
      POLYGON 31.800 25.300  31.800 26.300  32.800 26.300  32.800 25.300  
      31.800 25.300  ;
      POLYGON 31.800 23.300  31.800 24.300  32.800 24.300  32.800 23.300  
      31.800 23.300  ;
      POLYGON 31.800 21.300  31.800 22.300  32.800 22.300  32.800 21.300  
      31.800 21.300  ;
      POLYGON 29.300 3.200  29.300 4.200  30.300 4.200  30.300 3.200  29.300 
      3.200  ;
      POLYGON 26.800 23.300  26.800 24.300  27.800 24.300  27.800 23.300  
      26.800 23.300  ;
      POLYGON 26.800 25.300  26.800 26.300  27.800 26.300  27.800 25.300  
      26.800 25.300  ;
      POLYGON 25.800 3.200  25.800 4.200  26.800 4.200  26.800 3.200  25.800 
      3.200  ;
      POLYGON 23.800 25.300  23.800 26.300  24.800 26.300  24.800 25.300  
      23.800 25.300  ;
      POLYGON 23.800 23.300  23.800 24.300  24.800 24.300  24.800 23.300  
      23.800 23.300  ;
      POLYGON 23.800 21.300  23.800 22.300  24.800 22.300  24.800 21.300  
      23.800 21.300  ;
      POLYGON 20.800 3.200  20.800 4.200  21.800 4.200  21.800 3.200  20.800 
      3.200  ;
      POLYGON 20.800 25.300  20.800 26.300  21.800 26.300  21.800 25.300  
      20.800 25.300  ;
      POLYGON 20.800 23.300  20.800 24.300  21.800 24.300  21.800 23.300  
      20.800 23.300  ;
      POLYGON 20.800 21.300  20.800 22.300  21.800 22.300  21.800 21.300  
      20.800 21.300  ;
      POLYGON 15.800 3.200  15.800 4.200  16.800 4.200  16.800 3.200  15.800 
      3.200  ;
      POLYGON 15.800 23.300  15.800 24.300  16.800 24.300  16.800 23.300  
      15.800 23.300  ;
      POLYGON 15.800 25.300  15.800 26.300  16.800 26.300  16.800 25.300  
      15.800 25.300  ;
      POLYGON 15.800 21.300  15.800 22.300  16.800 22.300  16.800 21.300  
      15.800 21.300  ;
      POLYGON 10.800 3.200  10.800 4.200  11.800 4.200  11.800 3.200  10.800 
      3.200  ;
      POLYGON 10.800 25.300  10.800 26.300  11.800 26.300  11.800 25.300  
      10.800 25.300  ;
      POLYGON 10.800 23.300  10.800 24.300  11.800 24.300  11.800 23.300  
      10.800 23.300  ;
      POLYGON 10.800 21.300  10.800 22.300  11.800 22.300  11.800 21.300  
      10.800 21.300  ;
      POLYGON 7.300 3.200  7.300 4.200  8.300 4.200  8.300 3.200  7.300 3.200  ;
      
      POLYGON 7.300 21.300  7.300 22.300  8.300 22.300  8.300 21.300  7.300 
      21.300  ;
      POLYGON 7.300 23.300  7.300 24.300  8.300 24.300  8.300 23.300  7.300 
      23.300  ;
      POLYGON 7.300 25.300  7.300 26.300  8.300 26.300  8.300 25.300  7.300 
      25.300  ;
      POLYGON 4.300 3.200  4.300 4.200  5.300 4.200  5.300 3.200  4.300 3.200  ;
      
      POLYGON 4.300 25.300  4.300 26.300  5.300 26.300  5.300 25.300  4.300 
      25.300  ;
      POLYGON 4.300 21.300  4.300 22.300  5.300 22.300  5.300 21.300  4.300 
      21.300  ;
      POLYGON 4.300 23.300  4.300 24.300  5.300 24.300  5.300 23.300  4.300 
      23.300  ;
      POLYGON 1.300 25.300  1.300 26.300  2.300 26.300  2.300 25.300  1.300 
      25.300  ;
      POLYGON 1.300 3.200  1.300 4.200  2.300 4.200  2.300 3.200  1.300 3.200  ;
      
      POLYGON 1.300 21.300  1.300 22.300  2.300 22.300  2.300 21.300  1.300 
      21.300  ;
      POLYGON 1.300 23.300  1.300 24.300  2.300 24.300  2.300 23.300  1.300 
      23.300  ;
    LAYER FRAME ;
      POLYGON 0.000 0.000  56.000 0.000  56.000 30.000  0.000 30.000  0.000 
      0.000  ;
      RECT -0.500 28.500  56.500 30.500  ;
      RECT -0.500 -0.500  56.500 1.500  ;
    LAYER ML1 ;
      POLYGON 53.300 2.700  55.300 2.700  55.300 4.700  53.300 4.700  53.300 
      2.700  ;
      WIDTH 1.400  ;
      PATH 54.300 22.600 54.300 25.800  ;
      POLYGON 3.500 9.000  3.500 11.000  5.500 11.000  5.500 9.000  3.500 
      9.000  ;
      POLYGON 11.000 9.000  11.000 11.000  13.000 11.000  13.000 9.000  11.000 
      9.000  ;
      POLYGON 43.000 10.500  43.000 12.500  45.000 12.500  45.000 10.500  
      43.000 10.500  ;
      POLYGON 39.800 5.700  39.800 7.700  41.800 7.700  41.800 5.700  39.800 
      5.700  ;
      RECT 9.200 -0.500  11.200 1.500  ;
      RECT 26.700 -0.500  28.700 1.500  ;
      RECT 49.000 -0.500  51.000 1.500  ;
      RECT 37.300 17.700  39.300 19.700  ;
      RECT 37.300 13.000  39.300 15.000  ;
      RECT 30.300 15.700  32.300 17.700  ;
      RECT 27.300 17.700  29.300 19.700  ;
      RECT 21.300 9.000  23.300 11.000  ;
      RECT 21.300 17.700  23.300 19.700  ;
      RECT 16.300 15.000  18.300 17.000  ;
      RECT 11.000 9.000  13.000 11.000  ;
      RECT 3.500 9.000  5.500 11.000  ;
      RECT 9.200 28.500  11.200 30.500  ;
      RECT 26.700 28.500  28.700 30.500  ;
      RECT 49.000 28.500  51.000 30.500  ;
      RECT 53.300 24.800  55.300 26.800  ;
      RECT 53.300 22.800  55.300 24.800  ;
      RECT 53.300 20.800  55.300 22.800  ;
      RECT 53.300 2.700  55.300 4.700  ;
      RECT 50.300 24.800  52.300 26.800  ;
      RECT 50.300 22.800  52.300 24.800  ;
      RECT 50.300 20.800  52.300 22.800  ;
      RECT 50.300 2.700  52.300 4.700  ;
      RECT 47.300 24.800  49.300 26.800  ;
      RECT 47.300 22.800  49.300 24.800  ;
      RECT 47.300 20.800  49.300 22.800  ;
      RECT 47.300 2.700  49.300 4.700  ;
      RECT 43.800 2.700  45.800 4.700  ;
      RECT 42.300 20.800  44.300 22.800  ;
      RECT 42.300 22.800  44.300 24.800  ;
      RECT 42.300 24.800  44.300 26.800  ;
      RECT 39.300 24.800  41.300 26.800  ;
      RECT 39.300 22.800  41.300 24.800  ;
      RECT 39.300 20.800  41.300 22.800  ;
      RECT 38.800 2.700  40.800 4.700  ;
      RECT 36.300 24.800  38.300 26.800  ;
      RECT 36.300 22.800  38.300 24.800  ;
      RECT 36.300 20.800  38.300 22.800  ;
      RECT 33.800 2.700  35.800 4.700  ;
      RECT 31.300 24.800  33.300 26.800  ;
      RECT 31.300 22.800  33.300 24.800  ;
      RECT 31.300 20.800  33.300 22.800  ;
      RECT 28.800 2.700  30.800 4.700  ;
      RECT 26.300 22.800  28.300 24.800  ;
      RECT 26.300 24.800  28.300 26.800  ;
      RECT 25.300 2.700  27.300 4.700  ;
      RECT 23.300 24.800  25.300 26.800  ;
      RECT 23.300 22.800  25.300 24.800  ;
      RECT 23.300 20.800  25.300 22.800  ;
      RECT 20.300 2.700  22.300 4.700  ;
      RECT 20.300 24.800  22.300 26.800  ;
      RECT 20.300 22.800  22.300 24.800  ;
      RECT 20.300 20.800  22.300 22.800  ;
      RECT 15.300 2.700  17.300 4.700  ;
      RECT 15.300 22.800  17.300 24.800  ;
      RECT 15.300 24.800  17.300 26.800  ;
      RECT 15.300 20.800  17.300 22.800  ;
      RECT 10.300 2.700  12.300 4.700  ;
      RECT 10.300 24.800  12.300 26.800  ;
      RECT 10.300 22.800  12.300 24.800  ;
      RECT 10.300 20.800  12.300 22.800  ;
      RECT 6.800 2.700  8.800 4.700  ;
      RECT 6.800 20.800  8.800 22.800  ;
      RECT 6.800 22.800  8.800 24.800  ;
      RECT 6.800 24.800  8.800 26.800  ;
      RECT 3.800 2.700  5.800 4.700  ;
      RECT 3.800 24.800  5.800 26.800  ;
      RECT 3.800 20.800  5.800 22.800  ;
      RECT 3.800 22.800  5.800 24.800  ;
      RECT 0.800 24.800  2.800 26.800  ;
      RECT 0.800 2.700  2.800 4.700  ;
      RECT 0.800 20.800  2.800 22.800  ;
      RECT 0.800 22.800  2.800 24.800  ;
      POLYGON -0.500 30.500  -0.500 28.500  4.100 28.500  4.100 21.900  5.500 
      21.900  5.500 28.500  10.600 28.500  10.600 21.900  12.000 21.900  
      12.000 28.500  20.600 28.500  20.600 21.900  22.000 21.900  22.000 
      28.500  26.600 28.500  26.600 23.100  28.000 23.100  28.000 28.500  
      36.600 28.500  36.600 21.900  38.000 21.900  38.000 28.500  42.600 
      28.500  42.600 21.900  44.000 21.900  44.000 28.500  50.600 28.500  
      50.600 21.900  52.000 21.900  52.000 28.500  56.500 28.500  56.500 
      30.500  -0.500 30.500  ;
      POLYGON -0.500 1.500  -0.500 -0.500  56.500 -0.500  56.500 1.500  52.000 
      1.500  52.000 4.400  50.600 4.400  50.600 1.500  40.500 1.500  40.500 
      4.400  39.100 4.400  39.100 1.500  30.500 1.500  30.500 4.400  29.100 
      4.400  29.100 1.500  22.000 1.500  22.000 4.400  20.600 4.400  20.600 
      1.500  12.000 1.500  12.000 4.400  10.600 4.400  10.600 1.500  5.500 
      1.500  5.500 4.400  4.100 4.400  4.100 1.500  -0.500 1.500  ;
      POLYGON 1.100 26.500  1.100 21.900  1.300 21.900  1.300 3.000  2.300 
      3.000  2.300 6.200  4.800 6.200  4.800 5.700  6.800 5.700  6.800 7.700  
      4.800 7.700  4.800 7.200  2.300 7.200  2.300 12.500  4.300 12.500  4.300 
      12.000  6.300 12.000  6.300 14.000  4.300 14.000  4.300 13.500  2.300 
      13.500  2.300 18.300  4.800 18.300  4.800 17.800  6.800 17.800  6.800 
      19.800  4.800 19.800  4.800 19.300  2.300 19.300  2.300 21.900  2.500 
      21.900  2.500 26.500  1.100 26.500  ;
      POLYGON 7.300 16.700  7.300 9.000  7.800 9.000  7.800 3.000  8.800 3.000 
       8.800 6.200  13.800 6.200  13.800 5.700  15.800 5.700  15.800 7.700  
      13.800 7.700  13.800 7.200  8.800 7.200  8.800 10.000  8.300 10.000  
      8.300 15.700  31.800 15.700  31.800 16.700  8.800 16.700  8.800 26.500  
      7.800 26.500  7.800 16.700  7.300 16.700  ;
      POLYGON 9.300 14.000  9.300 12.000  11.300 12.000  11.300 12.500  14.300 
      12.500  14.300 12.000  16.300 12.000  16.300 12.500  27.300 12.500  
      27.300 12.000  29.300 12.000  29.300 12.500  34.000 12.500  34.000 
      12.700  34.300 12.700  34.300 14.700  32.300 14.700  32.300 13.500  
      29.300 13.500  29.300 14.000  27.300 14.000  27.300 13.500  16.300 
      13.500  16.300 14.000  14.300 14.000  14.300 13.500  11.300 13.500  
      11.300 14.000  9.300 14.000  ;
      POLYGON 15.800 4.700  15.800 3.200  16.800 3.200  16.800 3.700  17.300 
      3.700  17.300 9.500  21.300 9.500  21.300 9.000  23.300 9.000  23.300 
      11.000  21.300 11.000  21.300 10.500  16.300 10.500  16.300 4.700  
      15.800 4.700  ;
      POLYGON 15.600 26.500  15.600 21.900  15.800 21.900  15.800 18.300  
      21.300 18.300  21.300 17.700  23.300 17.700  23.300 19.700  21.300 
      19.700  21.300 19.300  16.800 19.300  16.800 21.900  17.000 21.900  
      17.000 26.500  15.600 26.500  ;
      POLYGON 19.300 7.700  19.300 5.700  21.300 5.700  21.300 6.200  25.600 
      6.200  25.600 2.700  27.000 2.700  27.000 5.700  28.300 5.700  28.300 
      7.700  26.300 7.700  26.300 7.200  21.300 7.200  21.300 7.700  19.300 
      7.700  ;
      POLYGON 24.300 11.000  24.300 9.000  26.300 9.000  26.300 9.700  44.300 
      9.700  44.300 10.500  45.000 10.500  45.000 12.500  43.000 12.500  
      43.000 10.700  26.300 10.700  26.300 11.000  24.300 11.000  ;
      POLYGON 26.300 7.700  26.300 5.700  28.300 5.700  28.300 7.700  26.300 
      7.700  ;
      POLYGON 23.600 26.500  23.600 21.100  23.800 21.100  23.800 20.800  
      27.300 20.800  27.300 17.700  29.300 17.700  29.300 19.700  28.300 
      19.700  28.300 21.800  25.000 21.800  25.000 26.500  23.600 26.500  ;
      POLYGON 31.600 26.500  31.600 21.900  31.800 21.900  31.800 18.700  
      37.300 18.700  37.300 17.700  39.300 17.700  39.300 19.700  32.800 
      19.700  32.800 21.900  33.000 21.900  33.000 26.500  31.600 26.500  ;
      POLYGON 34.300 7.200  34.300 3.200  35.300 3.200  35.300 6.200  39.800 
      6.200  39.800 5.700  41.800 5.700  41.800 7.700  39.800 7.700  39.800 
      7.200  34.300 7.200  ;
      POLYGON 44.800 8.700  44.800 3.200  45.800 3.200  45.800 7.700  50.300 
      7.700  50.300 9.700  49.000 9.700  49.000 14.500  41.300 14.500  41.300 
      16.700  48.300 16.700  48.300 16.200  50.300 16.200  50.300 18.200  
      48.300 18.200  48.300 17.700  41.300 17.700  41.300 22.000  41.000 
      22.000  41.000 26.500  39.600 26.500  39.600 21.900  40.300 21.900  
      40.300 14.500  37.900 14.500  37.900 13.500  48.000 13.500  48.000 8.700 
       44.800 8.700  ;
      POLYGON 47.800 6.700  47.800 3.000  48.800 3.000  48.800 5.700  53.300 
      5.700  53.300 7.700  52.500 7.700  52.500 17.900  53.300 17.900  53.300 
      19.900  48.700 19.900  48.700 21.900  49.000 21.900  49.000 26.500  
      47.600 26.500  47.600 21.900  47.700 21.900  47.700 18.900  51.300 
      18.900  51.300 17.900  51.500 17.900  51.500 7.700  51.300 7.700  51.300 
      6.700  47.800 6.700  ;
      POLYGON 53.500 12.500  53.500 10.500  54.300 10.500  54.300 2.700  
      55.300 2.700  55.300 10.500  55.500 10.500  55.500 12.500  55.300 12.500 
       55.300 26.500  54.300 26.500  54.300 12.500  53.500 12.500  ;
    LAYER ML2 ;
      POLYGON 3.500 9.000  3.500 11.000  5.500 11.000  5.500 9.000  3.500 
      9.000  ;
      POLYGON 11.000 11.000  11.000 9.000  13.000 9.000  13.000 11.000  11.000 
      11.000  ;
      POLYGON 21.300 11.000  21.300 9.000  23.300 9.000  23.300 11.000  22.800 
      11.000  22.800 17.700  23.300 17.700  23.300 19.700  21.300 19.700  
      21.300 17.700  21.800 17.700  21.800 11.000  21.300 11.000  ;
      POLYGON 26.300 7.700  26.300 5.700  28.300 5.700  28.300 6.200  28.800 
      6.200  28.800 17.700  29.300 17.700  29.300 19.700  27.300 19.700  
      27.300 17.700  27.800 17.700  27.800 7.700  26.300 7.700  ;
      POLYGON 37.300 19.700  37.300 17.700  37.800 17.700  37.800 7.200  
      39.800 7.200  39.800 5.700  41.800 5.700  41.800 7.700  41.300 7.700  
      41.300 8.200  38.800 8.200  38.800 17.700  39.300 17.700  39.300 19.700  
      37.300 19.700  ;
      POLYGON 43.000 12.500  43.000 10.500  45.000 10.500  45.000 12.500  
      43.000 12.500  ;
      POLYGON 53.500 12.500  53.500 10.500  55.500 10.500  55.500 12.500  
      53.500 12.500  ;
    LAYER POL ;
      POLYGON 2.800 27.800  2.800 1.700  3.800 1.700  3.800 9.000  5.500 9.000 
       5.500 11.000  3.800 11.000  3.800 27.800  2.800 27.800  ;
      POLYGON 4.800 19.800  4.800 17.800  6.800 17.800  6.800 27.800  5.800 
      27.800  5.800 19.800  4.800 19.800  ;
      POLYGON 4.300 14.000  4.300 12.000  6.300 12.000  6.300 12.500  9.300 
      12.500  9.300 12.000  11.300 12.000  11.300 14.000  9.300 14.000  9.300 
      13.500  6.300 13.500  6.300 14.000  4.300 14.000  ;
      POLYGON 4.800 7.700  4.800 5.700  5.800 5.700  5.800 1.700  6.800 1.700  
      6.800 7.700  4.800 7.700  ;
      POLYGON 11.000 11.000  11.000 9.000  12.300 9.000  12.300 1.900  13.300 
      1.900  13.300 27.600  12.300 27.600  12.300 11.000  11.000 11.000  ;
      POLYGON 13.800 7.700  13.800 5.700  14.300 5.700  14.300 1.900  15.300 
      1.900  15.300 5.700  15.800 5.700  15.800 7.700  13.800 7.700  ;
      POLYGON 14.300 27.600  14.300 11.000  17.300 11.000  17.300 1.900  
      18.300 1.900  18.300 12.000  16.300 12.000  16.300 14.000  15.300 14.000 
       15.300 27.600  14.300 27.600  ;
      POLYGON 16.300 17.000  16.300 15.000  18.300 15.000  18.300 27.600  
      17.300 27.600  17.300 17.000  16.300 17.000  ;
      POLYGON 19.300 27.500  19.300 1.800  20.300 1.800  20.300 5.700  21.300 
      5.700  21.300 7.700  20.300 7.700  20.300 27.500  19.300 27.500  ;
      POLYGON 21.300 19.700  21.300 17.700  23.300 17.700  23.300 27.600  
      22.300 27.600  22.300 19.700  21.300 19.700  ;
      POLYGON 21.300 11.000  21.300 9.000  22.300 9.000  22.300 1.900  23.300 
      1.900  23.300 11.000  21.300 11.000  ;
      POLYGON 24.300 15.000  24.300 1.900  25.300 1.900  25.300 9.000  26.300 
      9.000  26.300 11.000  25.300 11.000  25.300 14.000  26.300 14.000  
      26.300 27.600  25.300 27.600  25.300 15.000  24.300 15.000  ;
      POLYGON 26.300 7.700  26.300 5.700  26.800 5.700  26.800 5.200  30.800 
      5.200  30.800 1.900  31.800 1.900  31.800 6.200  28.300 6.200  28.300 
      7.700  26.300 7.700  ;
      POLYGON 27.300 14.000  27.300 12.000  27.800 12.000  27.800 8.700  
      29.500 8.700  29.500 7.200  32.800 7.200  32.800 1.900  33.800 1.900  
      33.800 8.200  30.500 8.200  30.500 9.700  28.800 9.700  28.800 12.000  
      29.300 12.000  29.300 14.000  27.300 14.000  ;
      POLYGON 30.300 27.600  30.300 10.700  35.800 10.700  35.800 1.900  
      36.800 1.900  36.800 11.700  31.300 11.700  31.300 15.700  32.300 15.700 
       32.300 17.700  31.300 17.700  31.300 27.600  30.300 27.600  ;
      POLYGON 27.300 19.700  27.300 17.700  29.300 17.700  29.300 27.600  
      28.300 27.600  28.300 19.700  27.300 19.700  ;
      POLYGON 32.300 14.700  32.300 12.700  34.300 12.700  34.300 27.600  
      33.300 27.600  33.300 14.700  32.300 14.700  ;
      POLYGON 35.300 27.600  35.300 13.500  37.300 13.500  37.300 13.000  
      37.800 13.000  37.800 1.900  38.800 1.900  38.800 13.000  39.300 13.000  
      39.300 15.000  37.300 15.000  37.300 14.500  36.300 14.500  36.300 
      27.600  35.300 27.600  ;
      POLYGON 39.800 7.700  39.800 5.700  40.800 5.700  40.800 1.900  41.800 
      1.900  41.800 7.700  39.800 7.700  ;
      POLYGON 41.300 27.600  41.300 11.500  42.800 11.500  42.800 1.900  
      43.800 1.900  43.800 10.500  45.000 10.500  45.000 12.500  42.300 12.500 
       42.300 27.600  41.300 27.600  ;
      POLYGON 37.300 19.700  37.300 17.700  39.300 17.700  39.300 27.600  
      38.300 27.600  38.300 19.700  37.300 19.700  ;
      POLYGON 48.300 9.700  48.300 7.700  49.300 7.700  49.300 1.900  50.300 
      1.900  50.300 9.700  48.300 9.700  ;
      POLYGON 51.300 7.700  51.300 5.700  52.300 5.700  52.300 1.900  53.300 
      1.900  53.300 7.700  51.300 7.700  ;
      POLYGON 48.300 18.200  48.300 16.200  50.300 16.200  50.300 27.600  
      49.300 27.600  49.300 18.200  48.300 18.200  ;
      POLYGON 51.300 19.900  51.300 17.900  53.300 17.900  53.300 27.600  
      52.300 27.600  52.300 19.900  51.300 19.900  ;
    LAYER VIA1 ;
      POLYGON 37.800 18.200  37.800 19.200  38.800 19.200  38.800 18.200  
      37.800 18.200  ;
      POLYGON 40.300 6.200  40.300 7.200  41.300 7.200  41.300 6.200  40.300 
      6.200  ;
      POLYGON 27.800 18.200  27.800 19.200  28.800 19.200  28.800 18.200  
      27.800 18.200  ;
      POLYGON 26.800 6.200  26.800 7.200  27.800 7.200  27.800 6.200  26.800 
      6.200  ;
      POLYGON 21.800 9.500  21.800 10.500  22.800 10.500  22.800 9.500  21.800 
      9.500  ;
      POLYGON 21.800 18.200  21.800 19.200  22.800 19.200  22.800 18.200  
      21.800 18.200  ;
      POLYGON 43.500 11.000  43.500 12.000  44.500 12.000  44.500 11.000  
      43.500 11.000  ;
      POLYGON 11.500 9.500  11.500 10.500  12.500 10.500  12.500 9.500  11.500 
      9.500  ;
      POLYGON 4.000 9.500  4.000 10.500  5.000 10.500  5.000 9.500  4.000 
      9.500  ;
      POLYGON 54.000 11.000  54.000 12.000  55.000 12.000  55.000 11.000  
      54.000 11.000  ;
  END
END sff1m2LEF


END LIBRARY
