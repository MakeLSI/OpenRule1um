*******************************************************************************
* CDL netlist
*
* Library : OpenRule1um
* Top Cell Name: rff1_r
* View Name: extracted
* Netlist created: 07.4.2020 15:03:09
*******************************************************************************

*.SCALE METER
*.GLOBAL vdd gnd

*******************************************************************************
* Library Name: OpenRule1um
* Cell Name:    rff1_r
* View Name:    extracted
*******************************************************************************

.SUBCKT rff1_r

MM88 n1 n9 n22 n2 pch w=6e-06 l=1e-06 as=3e-12 ps=8e-06 ad=6e-12 pd=1e-05 $X=4.23e-05 $Y=2.08e-05
MM86 n2 n3 n21 n2 pch w=6e-06 l=1e-06 as=6e-12 ps=8e-06 ad=1.2e-11 pd=1e-05 $X=3.73e-05 $Y=2.08e-05
MM66 n15 n3 n0 n0 nch w=2e-06 l=1e-06 as=2e-12 ps=6e-06 ad=1e-12 pd=4e-06 $X=2.58e-05 $Y=2.8e-06
MM84 n2 n7 n20 n2 pch w=6e-06 l=1e-06 as=3e-12 ps=8e-06 ad=6e-12 pd=1e-05 $X=2.88e-05 $Y=2.08e-05
MM90 n2 n1 n23 n2 pch w=6e-06 l=1e-06 as=3e-12 ps=8e-06 ad=6e-12 pd=1e-05 $X=4.73e-05 $Y=2.08e-05
MM60 n0 n13 n12 n0 nch w=2e-06 l=1e-06 as=4e-12 ps=6e-06 ad=4e-12 pd=6e-06 $X=2.8e-06 $Y=2.8e-06
MM82 n7 n8 n19 n2 pch w=6e-06 l=1e-06 as=3e-12 ps=8e-06 ad=6e-12 pd=1e-05 $X=2.38e-05 $Y=2.08e-05
MM87 n21 n8 n1 n2 pch w=6e-06 l=1e-06 as=6e-12 ps=1e-05 ad=3e-12 pd=8e-06 $X=3.93e-05 $Y=2.08e-05
MM91 n23 n6 n4 n2 pch w=6e-06 l=1e-06 as=6e-12 ps=1e-05 ad=3e-12 pd=8e-06 $X=4.93e-05 $Y=2.08e-05
MM78 n9 n12 n2 n2 pch w=6e-06 l=1e-06 as=1.2e-11 ps=1e-05 ad=1.2e-11 pd=1e-05 $X=9.3e-06 $Y=2.08e-05
MM71 n1 n8 n17 n0 nch w=2e-06 l=1e-06 as=1e-12 ps=4e-06 ad=2e-12 pd=6e-06 $X=3.98e-05 $Y=2.8e-06
MM73 n0 n1 n4 n0 nch w=2e-06 l=1e-06 as=2e-12 ps=6e-06 ad=2e-12 pd=6e-06 $X=4.48e-05 $Y=2.8e-06
MM77 n2 n13 n12 n2 pch w=6e-06 l=1e-06 as=1.2e-11 ps=1e-05 ad=1.2e-11 pd=1e-05 $X=2.8e-06 $Y=1.95e-05
MM61 n9 n12 n0 n0 nch w=2e-06 l=1e-06 as=4e-12 ps=6e-06 ad=4e-12 pd=6e-06 $X=9.3e-06 $Y=2.8e-06
MM75 n5 n4 n0 n0 nch w=2e-06 l=1e-06 as=4e-12 ps=6e-06 ad=4e-12 pd=6e-06 $X=5.58e-05 $Y=2.8e-06
MM92 n5 n4 n2 n2 pch w=6e-06 l=1e-06 as=1.2e-11 ps=1e-05 ad=1.2e-11 pd=1e-05 $X=5.58e-05 $Y=2.08e-05
MM74 n4 n6 n0 n0 nch w=2e-06 l=1e-06 as=1.9e-12 ps=5.8e-06 ad=2e-12 pd=6e-06 $X=4.78e-05 $Y=2.8e-06
MM79 n2 n9 n8 n2 pch w=6e-06 l=1e-06 as=6e-12 ps=1e-05 ad=6e-12 pd=1e-05 $X=1.23e-05 $Y=2.08e-05
MM69 n0 n3 n16 n0 nch w=2e-06 l=1e-06 as=1e-12 ps=4e-06 ad=2e-12 pd=6e-06 $X=3.48e-05 $Y=2.8e-06
MM63 n0 n10 n14 n0 nch w=2e-06 l=1e-06 as=2e-12 ps=4e-06 ad=4e-12 pd=6e-06 $X=1.88e-05 $Y=2.8e-06
MM67 n0 n7 n3 n0 nch w=2e-06 l=1e-06 as=2e-12 ps=6e-06 ad=2e-12 pd=6e-06 $X=2.88e-05 $Y=2.8e-06
MM83 n19 n3 n2 n2 pch w=6e-06 l=1e-06 as=6e-12 ps=1e-05 ad=3e-12 pd=8e-06 $X=2.58e-05 $Y=2.08e-05
MM65 n7 n9 n15 n0 nch w=2e-06 l=1e-06 as=1e-12 ps=4e-06 ad=2e-12 pd=6e-06 $X=2.38e-05 $Y=2.8e-06
MM80 n2 n10 n18 n2 pch w=6e-06 l=1e-06 as=6e-12 ps=8e-06 ad=1.2e-11 pd=1e-05 $X=1.88e-05 $Y=2.08e-05
MM62 n0 n9 n8 n0 nch w=2e-06 l=1e-06 as=2e-12 ps=6e-06 ad=2e-12 pd=6e-06 $X=1.23e-05 $Y=2.8e-06
MM76 n0 n5 n11 n0 nch w=2e-06 l=1e-06 as=2e-12 ps=6e-06 ad=2e-12 pd=6e-06 $X=5.88e-05 $Y=2.8e-06
MM89 n22 n4 n2 n2 pch w=6e-06 l=1e-06 as=6e-12 ps=1e-05 ad=3e-12 pd=8e-06 $X=4.43e-05 $Y=2.08e-05
MM70 n16 n9 n1 n0 nch w=2e-06 l=1e-06 as=2e-12 ps=6e-06 ad=1e-12 pd=4e-06 $X=3.68e-05 $Y=2.8e-06
MM81 n18 n9 n7 n2 pch w=6e-06 l=1e-06 as=6e-12 ps=1e-05 ad=3e-12 pd=8e-06 $X=2.08e-05 $Y=2.08e-05
MM85 n20 n6 n3 n2 pch w=6e-06 l=1e-06 as=6e-12 ps=1e-05 ad=3e-12 pd=8e-06 $X=3.08e-05 $Y=2.08e-05
MM68 n3 n6 n0 n0 nch w=2e-06 l=1e-06 as=2e-12 ps=6e-06 ad=2e-12 pd=6e-06 $X=3.18e-05 $Y=2.8e-06
MM93 n2 n5 n11 n2 pch w=6e-06 l=1e-06 as=6e-12 ps=1e-05 ad=6e-12 pd=1e-05 $X=5.88e-05 $Y=2.08e-05
MM64 n14 n8 n7 n0 nch w=2e-06 l=1e-06 as=2e-12 ps=6e-06 ad=1e-12 pd=4e-06 $X=2.08e-05 $Y=2.8e-06
MM72 n17 n4 n0 n0 nch w=2e-06 l=1e-06 as=2e-12 ps=6e-06 ad=1e-12 pd=4e-06 $X=4.18e-05 $Y=2.8e-06
.ENDS
