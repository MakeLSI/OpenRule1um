*******************************************************************************
* CDL netlist
*
* Library : OpenRule1um
* Top Cell Name: rff1_r
* View Name: schematic
* Netlist created: 07.4.2020 15:03:09
*******************************************************************************

*.SCALE METER
*.GLOBAL vdd gnd

*******************************************************************************
* Library Name: OpenRule1um
* Cell Name:    rff1_r
* View Name:    schematic
*******************************************************************************

.SUBCKT rff1_r CK S VDD Q D VSS 
*.PININFO CK:I VDD:B S:I Q:O D:I VSS:B QB:O

M29 n4 n25 VSS VSS nch w=2u l=1u m=1
M2 n19 n17 n15 VDD pch w=6u l=1u m=1
M20 n25 n18 n24 VSS nch w=2u l=1u m=1
M24 n26 n18 n25 VDD pch w=6u l=1u m=1
M26 n25 n17 n9 VSS nch w=2u l=1u m=1
M27 n24 n4 VSS VSS nch w=2u l=1u m=1
M22 VDD n4 n8 VDD pch w=6u l=1u m=1
M0 VDD n17 n18 VDD pch w=6u l=1u m=1
M14 n5 S n22 VDD pch w=6u l=1u m=1
M12 VDD n15 n5 VDD pch w=6u l=1u m=1
M4 n15 n18 n20 VSS nch w=2u l=1u m=1
M6 n17 n2 VSS VSS nch w=2u l=1u m=1
M17 n28 S n4 VDD pch w=6u l=1u m=1
M23 n9 n22 VSS VSS nch w=2u l=1u m=1
M28 n4 S VSS VSS nch w=2u l=1u m=1
M19 VDD n25 n28 VDD pch w=6u l=1u m=1
M11 n15 n17 n14 VSS nch w=2u l=1u m=1
M16 n22 n15 VSS VSS nch w=2u l=1u m=1
M9 n14 n22 VSS VSS nch w=2u l=1u m=1
M34 n2 CK VSS VSS nch w=2u l=1u m=1
M15 n22 S VSS VSS nch w=2u l=1u m=1
M25 VDD n22 n26 VDD pch w=6u l=1u m=1
M30 VDD n4 QB VDD pch w=6u l=1u m=1
M5 n20 D VSS VSS nch w=2u l=1u m=1
M32_40 Q QB VSS VSS nch w=2u l=1u m=1
M3 VDD D n19 VDD pch w=6u l=1u m=1
M21 n8 n17 n25 VDD pch w=6u l=1u m=1
M32 VDD CK n2 VDD pch w=6u l=1u m=1
M8 VDD n22 n21 VDD pch w=6u l=1u m=1
M7 VDD n2 n17 VDD pch w=6u l=1u m=1
M31 VDD QB Q VDD pch w=6u l=1u m=1
M1 n18 n17 VSS VSS nch w=2u l=1u m=1
M33 QB n4 VSS VSS nch w=2u l=1u m=1
M10 n21 n18 n15 VDD pch w=6u l=1u m=1
.ENDS

