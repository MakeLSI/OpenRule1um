VERSION 5.3 ;

NAMESCASESENSITIVE ON ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS











MACRO inv1LEF
  CLASS BLOCK ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER POL ;
        POLYGON 1.000 16.500  1.000 14.500  2.800 14.500  2.800 1.700  3.800 
        1.700  3.800 26.500  2.800 26.500  2.800 16.500  1.000 16.500  ;
    END
    PORT
      LAYER ML1 ;
        RECT 1.000 14.500  3.000 16.500  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    PORT
      LAYER ML1 ;
        POLYGON -0.500 30.500  -0.500 28.500  1.100 28.500  1.100 20.600  
        2.500 20.600  2.500 28.500  7.000 28.500  7.000 30.500  -0.500 30.500  ;
        
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    PORT
      LAYER ML1 ;
        POLYGON -0.500 1.500  -0.500 -0.500  7.000 -0.500  7.000 1.500  2.300 
        1.500  2.300 4.200  1.300 4.200  1.300 1.500  -0.500 1.500  ;
    END
  END VSS
  PIN YB
    DIRECTION OUTPUT ;
    PORT
      LAYER ML1 ;
        POLYGON 4.000 12.300  4.000 10.300  4.300 10.300  4.300 3.200  5.300 
        3.200  5.300 10.300  6.000 10.300  6.000 12.300  5.300 12.300  5.300 
        20.600  5.500 20.600  5.500 25.200  4.100 25.200  4.100 20.600  4.300 
        20.600  4.300 12.300  4.000 12.300  ;
    END
  END YB
  OBS
    LAYER CNT ;
      POLYGON 1.300 22.000  1.300 23.000  2.300 23.000  2.300 22.000  1.300 
      22.000  ;
      POLYGON 1.300 20.000  1.300 21.000  2.300 21.000  2.300 20.000  1.300 
      20.000  ;
      POLYGON 1.300 3.200  1.300 4.200  2.300 4.200  2.300 3.200  1.300 3.200  ;
      
      POLYGON 1.300 24.000  1.300 25.000  2.300 25.000  2.300 24.000  1.300 
      24.000  ;
      POLYGON 4.300 22.000  4.300 23.000  5.300 23.000  5.300 22.000  4.300 
      22.000  ;
      POLYGON 4.300 20.000  4.300 21.000  5.300 21.000  5.300 20.000  4.300 
      20.000  ;
      POLYGON 4.300 24.000  4.300 25.000  5.300 25.000  5.300 24.000  4.300 
      24.000  ;
      POLYGON 4.300 3.200  4.300 4.200  5.300 4.200  5.300 3.200  4.300 3.200  ;
      
      POLYGON 3.000 29.000  3.000 30.000  4.000 30.000  4.000 29.000  3.000 
      29.000  ;
      POLYGON 1.500 15.000  1.500 16.000  2.500 16.000  2.500 15.000  1.500 
      15.000  ;
      POLYGON 3.500 0.000  3.500 1.000  4.500 1.000  4.500 0.000  3.500 0.000  ;
      
    LAYER FRAME ;
      POLYGON 0.000 0.000  6.500 0.000  6.500 30.000  0.000 30.000  0.000 
      0.000  ;
      RECT -0.500 -0.500  7.000 1.500  ;
      RECT -0.500 28.500  7.000 30.500  ;
    LAYER ML1 ;
      RECT 2.500 28.500  4.500 30.500  ;
      RECT 1.000 14.500  3.000 16.500  ;
      RECT 3.000 -0.500  5.000 1.500  ;
      POLYGON 1.000 14.500  1.000 16.500  3.000 16.500  3.000 14.500  1.000 
      14.500  ;
      RECT 3.800 2.700  5.800 4.700  ;
      RECT 3.800 23.500  5.800 25.500  ;
      RECT 3.800 19.500  5.800 21.500  ;
      RECT 3.800 21.500  5.800 23.500  ;
      RECT 0.800 23.500  2.800 25.500  ;
      RECT 0.800 2.700  2.800 4.700  ;
      RECT 0.800 19.500  2.800 21.500  ;
      RECT 0.800 21.500  2.800 23.500  ;
      POLYGON -0.500 30.500  -0.500 28.500  1.100 28.500  1.100 20.600  2.500 
      20.600  2.500 28.500  7.000 28.500  7.000 30.500  -0.500 30.500  ;
      POLYGON -0.500 1.500  -0.500 -0.500  7.000 -0.500  7.000 1.500  2.300 
      1.500  2.300 4.200  1.300 4.200  1.300 1.500  -0.500 1.500  ;
      POLYGON 4.000 12.300  4.000 10.300  4.300 10.300  4.300 3.200  5.300 
      3.200  5.300 10.300  6.000 10.300  6.000 12.300  5.300 12.300  5.300 
      20.600  5.500 20.600  5.500 25.200  4.100 25.200  4.100 20.600  4.300 
      20.600  4.300 12.300  4.000 12.300  ;
    LAYER ML2 ;
      POLYGON 4.000 10.300  4.000 12.300  6.000 12.300  6.000 10.300  4.000 
      10.300  ;
      POLYGON 1.000 14.500  1.000 16.500  3.000 16.500  3.000 14.500  1.000 
      14.500  ;
    LAYER POL ;
      POLYGON 1.000 16.500  1.000 14.500  2.800 14.500  2.800 1.700  3.800 
      1.700  3.800 26.500  2.800 26.500  2.800 16.500  1.000 16.500  ;
    LAYER VIA1 ;
      POLYGON 4.500 10.800  4.500 11.800  5.500 11.800  5.500 10.800  4.500 
      10.800  ;
      POLYGON 1.500 15.000  1.500 16.000  2.500 16.000  2.500 15.000  1.500 
      15.000  ;
  END
END inv1LEF


END LIBRARY
