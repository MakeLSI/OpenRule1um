VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO nr212
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 12.500 BY 30.000 ;
  SYMMETRY X Y ;
  SITE unit ;
 
  PIN A0
    USE SIGNAL ;
    PORT
      LAYER ML1 ;
        POLYGON 1.000 14.500  1.000 16.500  3.000 16.500  3.000 14.500  1.000 
        14.500  ;
    END
    PORT
      LAYER ML2 ;
        POLYGON 1.000 14.500  1.000 16.500  3.000 16.500  3.000 14.500  1.000 
        14.500  ;
    END
  END A0
  PIN A1
    USE SIGNAL ;
    PORT
      LAYER ML1 ;
        POLYGON 4.000 8.500  4.000 10.500  6.000 10.500  6.000 8.500  4.000 
        8.500  ;
    END
    PORT
      LAYER ML2 ;
        POLYGON 4.000 8.500  4.000 10.500  6.000 10.500  6.000 8.500  4.000 
        8.500  ;
    END
  END A1
  PIN B0
    USE SIGNAL ;
    PORT
      LAYER ML1 ;
        POLYGON 7.000 11.500  7.000 13.500  9.000 13.500  9.000 11.500  7.000 
        11.500  ;
    END
    PORT
      LAYER ML2 ;
        POLYGON 7.000 11.500  7.000 13.500  9.000 13.500  9.000 11.500  7.000 
        11.500  ;
    END
  END B0
  PIN VDD
    USE POWER ;
    PORT
      LAYER ML1 ;
        RECT -0.500 28.500  13.000 30.500  ;
    END
  END VDD
  PIN VSS
    USE GROUND ;
    PORT
      LAYER ML1 ;
        RECT -0.500 -0.500  13.000 1.500  ;
    END
  END VSS
  PIN YB
    USE SIGNAL ;
    PORT
      LAYER ML1 ;
        WIDTH 1.000  ;
        PATH 10.800 20.500 10.800 18.000 10.500 18.000 10.500 6.500 6.800 
        6.500 6.800 3.800  ;
    END
    PORT
      LAYER ML1 ;
        POLYGON 9.500 8.500  9.500 10.500  11.500 10.500  11.500 8.500  9.500 
        8.500  ;
    END
    PORT
      LAYER ML2 ;
        POLYGON 9.500 8.500  9.500 10.500  11.500 10.500  11.500 8.500  9.500 
        8.500  ;
    END
  END YB
  OBS

    LAYER ML1 ;

      WIDTH 1.000  ;
      PATH 1.800 24.500 1.800 18.000 7.800 18.000 7.800 24.500  ;
      WIDTH 1.000  ;
      PATH 10.800 20.500 10.800 18.000 10.500 18.000 10.500 6.500 6.800 6.500 
      6.800 3.800  ;
      WIDTH 1.400  ;
      PATH 10.800 21.300 10.800 24.500  ;

      WIDTH 1.000  ;
      PATH 9.800 1.000 9.800 3.800  ;
      WIDTH 1.400  ;
      PATH 4.800 21.300 4.800 28.500  ;
      WIDTH 1.000  ;
      PATH 1.800 1.000 1.800 3.800  ;
      WIDTH 1.400  ;
      PATH 1.800 21.300 1.800 24.500  ;

    VIA 1.800 22.500  dcont ;
    VIA 1.800 20.500  dcont ;
    VIA 1.800 3.800  dcont ;
    VIA 1.800 24.500  dcont ;
    VIA 4.800 22.500  dcont ;
    VIA 4.800 20.500  dcont ;
    VIA 4.800 24.500  dcont ;
    VIA 6.800 3.800  dcont ;
    VIA 7.800 24.500  dcont ;
    VIA 7.800 22.500  dcont ;
    VIA 7.800 20.500  dcont ;
    VIA 9.800 3.800  dcont ;
    VIA 10.800 20.500  dcont ;
    VIA 10.800 22.500  dcont ;
    VIA 10.800 24.500  dcont ;
    VIA 5.000 9.500  pcont ;
    VIA 7.000 29.500  nsubcont ;
    VIA 8.000 12.500  pcont ;
    VIA 2.000 15.500  pcont ;
    VIA 6.000 0.500  psubcont ;
  END
END nr212

MACRO dcont
  CLASS CORE ;
  OBS
    LAYER ML1 ;
      RECT -1.000 -1.000  1.000 1.000  ;
  END
END dcont

MACRO pcont
  CLASS CORE ;
  OBS
    LAYER ML1 ;
      RECT -1.000 -1.000  1.000 1.000  ;
  END
END pcont

MACRO nsubcont
  CLASS CORE ;
  OBS
    LAYER ML1 ;
      RECT -1.000 -1.000  1.000 1.000  ;
  END
END nsubcont

MACRO psubcont
  CLASS CORE ;
  OBS
    LAYER ML1 ;
      RECT -1.000 -1.000  1.000 1.000  ;
  END
END psubcont


END LIBRARY
