VERSION 5.3 ;

NAMESCASESENSITIVE ON ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS











MACRO inv8LEF
  CLASS BLOCK ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER POL ;
        POLYGON 1.000 16.500  1.000 14.500  2.800 14.500  2.800 1.700  3.800 
        1.700  3.800 14.500  5.800 14.500  5.800 1.700  6.800 1.700  6.800 
        14.500  8.800 14.500  8.800 1.700  9.800 1.700  9.800 14.500  11.800 
        14.500  11.800 1.700  12.800 1.700  12.800 14.500  14.800 14.500  
        14.800 1.700  15.800 1.700  15.800 14.500  17.800 14.500  17.800 1.700 
         18.800 1.700  18.800 14.500  20.800 14.500  20.800 1.700  21.800 
        1.700  21.800 14.500  23.800 14.500  23.800 1.700  24.800 1.700  
        24.800 26.500  23.800 26.500  23.800 16.500  21.800 16.500  21.800 
        26.500  20.800 26.500  20.800 16.500  18.800 16.500  18.800 26.500  
        17.800 26.500  17.800 16.500  15.800 16.500  15.800 26.500  14.800 
        26.500  14.800 16.500  12.800 16.500  12.800 26.500  11.800 26.500  
        11.800 16.500  9.800 16.500  9.800 26.500  8.800 26.500  8.800 16.500  
        6.800 16.500  6.800 26.500  5.800 26.500  5.800 16.500  3.800 16.500  
        3.800 26.500  2.800 26.500  2.800 16.500  1.000 16.500  ;
    END
    PORT
      LAYER ML1 ;
        POLYGON 1.000 14.500  1.000 16.500  3.000 16.500  3.000 14.500  1.000 
        14.500  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    PORT
      LAYER ML1 ;
        POLYGON -0.500 30.500  -0.500 28.500  1.100 28.500  1.100 20.600  
        2.500 20.600  2.500 28.500  7.100 28.500  7.100 20.600  8.500 20.600  
        8.500 28.500  13.100 28.500  13.100 20.600  14.500 20.600  14.500 
        28.500  19.100 28.500  19.100 20.600  20.500 20.600  20.500 28.500  
        25.100 28.500  25.100 20.600  26.500 20.600  26.500 28.500  28.000 
        28.500  28.000 30.500  -0.500 30.500  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    PORT
      LAYER ML1 ;
        POLYGON -0.500 1.500  -0.500 -0.500  28.000 -0.500  28.000 1.500  
        26.300 1.500  26.300 4.200  25.300 4.200  25.300 1.500  20.300 1.500  
        20.300 4.200  19.300 4.200  19.300 1.500  14.300 1.500  14.300 4.200  
        13.300 4.200  13.300 1.500  8.300 1.500  8.300 4.200  7.300 4.200  
        7.300 1.500  2.300 1.500  2.300 4.200  1.300 4.200  1.300 1.500  
        -0.500 1.500  ;
    END
  END VSS
  PIN YB
    DIRECTION OUTPUT ;
    PORT
      LAYER ML1 ;
        POLYGON 4.100 25.200  4.100 20.600  4.300 20.600  4.300 3.200  5.300 
        3.200  5.300 10.500  10.300 10.500  10.300 3.200  11.300 3.200  11.300 
        10.500  16.300 10.500  16.300 3.200  17.300 3.200  17.300 10.500  
        22.300 10.500  22.300 3.200  23.300 3.200  23.300 10.500  24.000 
        10.500  24.000 12.500  23.300 12.500  23.300 20.600  23.500 20.600  
        23.500 25.200  22.100 25.200  22.100 20.600  22.300 20.600  22.300 
        12.500  22.000 12.500  22.000 11.500  17.300 11.500  17.300 20.600  
        17.500 20.600  17.500 25.200  16.100 25.200  16.100 20.600  16.300 
        20.600  16.300 11.500  11.300 11.500  11.300 20.600  11.500 20.600  
        11.500 25.200  10.100 25.200  10.100 20.600  10.300 20.600  10.300 
        11.500  5.300 11.500  5.300 20.600  5.500 20.600  5.500 25.200  4.100 
        25.200  ;
    END
  END YB
  OBS
    LAYER CNT ;
      POLYGON 22.300 20.000  22.300 21.000  23.300 21.000  23.300 20.000  
      22.300 20.000  ;
      POLYGON 22.300 3.200  22.300 4.200  23.300 4.200  23.300 3.200  22.300 
      3.200  ;
      POLYGON 25.300 22.000  25.300 23.000  26.300 23.000  26.300 22.000  
      25.300 22.000  ;
      POLYGON 25.300 20.000  25.300 21.000  26.300 21.000  26.300 20.000  
      25.300 20.000  ;
      POLYGON 25.300 24.000  25.300 25.000  26.300 25.000  26.300 24.000  
      25.300 24.000  ;
      POLYGON 25.300 3.200  25.300 4.200  26.300 4.200  26.300 3.200  25.300 
      3.200  ;
      POLYGON 4.500 29.000  4.500 30.000  5.500 30.000  5.500 29.000  4.500 
      29.000  ;
      POLYGON 17.800 0.000  17.800 1.000  18.800 1.000  18.800 0.000  17.800 
      0.000  ;
      POLYGON 1.500 15.000  1.500 16.000  2.500 16.000  2.500 15.000  1.500 
      15.000  ;
      POLYGON 4.500 0.000  4.500 1.000  5.500 1.000  5.500 0.000  4.500 0.000  ;
      
      POLYGON 18.600 29.000  18.600 30.000  19.600 30.000  19.600 29.000  
      18.600 29.000  ;
      POLYGON 22.300 22.000  22.300 23.000  23.300 23.000  23.300 22.000  
      22.300 22.000  ;
      POLYGON 22.300 24.000  22.300 25.000  23.300 25.000  23.300 24.000  
      22.300 24.000  ;
      POLYGON 19.300 3.200  19.300 4.200  20.300 4.200  20.300 3.200  19.300 
      3.200  ;
      POLYGON 19.300 22.000  19.300 23.000  20.300 23.000  20.300 22.000  
      19.300 22.000  ;
      POLYGON 19.300 20.000  19.300 21.000  20.300 21.000  20.300 20.000  
      19.300 20.000  ;
      POLYGON 19.300 24.000  19.300 25.000  20.300 25.000  20.300 24.000  
      19.300 24.000  ;
      POLYGON 16.300 3.200  16.300 4.200  17.300 4.200  17.300 3.200  16.300 
      3.200  ;
      POLYGON 16.300 22.000  16.300 23.000  17.300 23.000  17.300 22.000  
      16.300 22.000  ;
      POLYGON 16.300 20.000  16.300 21.000  17.300 21.000  17.300 20.000  
      16.300 20.000  ;
      POLYGON 16.300 24.000  16.300 25.000  17.300 25.000  17.300 24.000  
      16.300 24.000  ;
      POLYGON 13.300 3.200  13.300 4.200  14.300 4.200  14.300 3.200  13.300 
      3.200  ;
      POLYGON 13.300 24.000  13.300 25.000  14.300 25.000  14.300 24.000  
      13.300 24.000  ;
      POLYGON 13.300 22.000  13.300 23.000  14.300 23.000  14.300 22.000  
      13.300 22.000  ;
      POLYGON 13.300 20.000  13.300 21.000  14.300 21.000  14.300 20.000  
      13.300 20.000  ;
      POLYGON 10.300 3.200  10.300 4.200  11.300 4.200  11.300 3.200  10.300 
      3.200  ;
      POLYGON 10.300 22.000  10.300 23.000  11.300 23.000  11.300 22.000  
      10.300 22.000  ;
      POLYGON 10.300 20.000  10.300 21.000  11.300 21.000  11.300 20.000  
      10.300 20.000  ;
      POLYGON 10.300 24.000  10.300 25.000  11.300 25.000  11.300 24.000  
      10.300 24.000  ;
      POLYGON 7.300 24.000  7.300 25.000  8.300 25.000  8.300 24.000  7.300 
      24.000  ;
      POLYGON 7.300 22.000  7.300 23.000  8.300 23.000  8.300 22.000  7.300 
      22.000  ;
      POLYGON 7.300 20.000  7.300 21.000  8.300 21.000  8.300 20.000  7.300 
      20.000  ;
      POLYGON 7.300 3.200  7.300 4.200  8.300 4.200  8.300 3.200  7.300 3.200  ;
      
      POLYGON 4.300 24.000  4.300 25.000  5.300 25.000  5.300 24.000  4.300 
      24.000  ;
      POLYGON 4.300 20.000  4.300 21.000  5.300 21.000  5.300 20.000  4.300 
      20.000  ;
      POLYGON 4.300 22.000  4.300 23.000  5.300 23.000  5.300 22.000  4.300 
      22.000  ;
      POLYGON 4.300 3.200  4.300 4.200  5.300 4.200  5.300 3.200  4.300 3.200  ;
      
      POLYGON 1.300 24.000  1.300 25.000  2.300 25.000  2.300 24.000  1.300 
      24.000  ;
      POLYGON 1.300 20.000  1.300 21.000  2.300 21.000  2.300 20.000  1.300 
      20.000  ;
      POLYGON 1.300 22.000  1.300 23.000  2.300 23.000  2.300 22.000  1.300 
      22.000  ;
      POLYGON 1.300 3.200  1.300 4.200  2.300 4.200  2.300 3.200  1.300 3.200  ;
      
    LAYER FRAME ;
      RECT -0.500 28.500  28.000 30.500  ;
      RECT -0.500 -0.500  28.000 1.500  ;
      POLYGON 0.000 0.000  27.500 0.000  27.500 30.000  0.000 30.000  0.000 
      0.000  ;
    LAYER ML1 ;
      WIDTH 1.400  ;
      PATH 19.800 21.300 19.800 24.500  ;
      WIDTH 1.400  ;
      PATH 25.800 21.300 25.800 24.500  ;
      POLYGON 1.000 14.500  1.000 16.500  3.000 16.500  3.000 14.500  1.000 
      14.500  ;
      RECT 18.100 28.500  20.100 30.500  ;
      RECT 4.000 -0.500  6.000 1.500  ;
      RECT 1.000 14.500  3.000 16.500  ;
      RECT 17.300 -0.500  19.300 1.500  ;
      RECT 4.000 28.500  6.000 30.500  ;
      RECT 24.800 2.700  26.800 4.700  ;
      RECT 24.800 23.500  26.800 25.500  ;
      RECT 24.800 19.500  26.800 21.500  ;
      RECT 24.800 21.500  26.800 23.500  ;
      RECT 21.800 2.700  23.800 4.700  ;
      RECT 21.800 19.500  23.800 21.500  ;
      RECT 21.800 21.500  23.800 23.500  ;
      RECT 21.800 23.500  23.800 25.500  ;
      RECT 18.800 2.700  20.800 4.700  ;
      RECT 18.800 21.500  20.800 23.500  ;
      RECT 18.800 19.500  20.800 21.500  ;
      RECT 18.800 23.500  20.800 25.500  ;
      RECT 15.800 2.700  17.800 4.700  ;
      RECT 15.800 21.500  17.800 23.500  ;
      RECT 15.800 19.500  17.800 21.500  ;
      RECT 15.800 23.500  17.800 25.500  ;
      RECT 12.800 2.700  14.800 4.700  ;
      RECT 12.800 23.500  14.800 25.500  ;
      RECT 12.800 21.500  14.800 23.500  ;
      RECT 12.800 19.500  14.800 21.500  ;
      RECT 9.800 2.700  11.800 4.700  ;
      RECT 9.800 21.500  11.800 23.500  ;
      RECT 9.800 19.500  11.800 21.500  ;
      RECT 9.800 23.500  11.800 25.500  ;
      RECT 6.800 23.500  8.800 25.500  ;
      RECT 6.800 21.500  8.800 23.500  ;
      RECT 6.800 19.500  8.800 21.500  ;
      RECT 6.800 2.700  8.800 4.700  ;
      RECT 3.800 23.500  5.800 25.500  ;
      RECT 3.800 19.500  5.800 21.500  ;
      RECT 3.800 21.500  5.800 23.500  ;
      RECT 3.800 2.700  5.800 4.700  ;
      RECT 0.800 23.500  2.800 25.500  ;
      RECT 0.800 19.500  2.800 21.500  ;
      RECT 0.800 21.500  2.800 23.500  ;
      RECT 0.800 2.700  2.800 4.700  ;
      POLYGON -0.500 30.500  -0.500 28.500  1.100 28.500  1.100 20.600  2.500 
      20.600  2.500 28.500  7.100 28.500  7.100 20.600  8.500 20.600  8.500 
      28.500  13.100 28.500  13.100 20.600  14.500 20.600  14.500 28.500  
      19.100 28.500  19.100 20.600  20.500 20.600  20.500 28.500  25.100 
      28.500  25.100 20.600  26.500 20.600  26.500 28.500  28.000 28.500  
      28.000 30.500  -0.500 30.500  ;
      POLYGON -0.500 1.500  -0.500 -0.500  28.000 -0.500  28.000 1.500  26.300 
      1.500  26.300 4.200  25.300 4.200  25.300 1.500  20.300 1.500  20.300 
      4.200  19.300 4.200  19.300 1.500  14.300 1.500  14.300 4.200  13.300 
      4.200  13.300 1.500  8.300 1.500  8.300 4.200  7.300 4.200  7.300 1.500  
      2.300 1.500  2.300 4.200  1.300 4.200  1.300 1.500  -0.500 1.500  ;
      POLYGON 4.100 25.200  4.100 20.600  4.300 20.600  4.300 3.200  5.300 
      3.200  5.300 10.500  10.300 10.500  10.300 3.200  11.300 3.200  11.300 
      10.500  16.300 10.500  16.300 3.200  17.300 3.200  17.300 10.500  22.300 
      10.500  22.300 3.200  23.300 3.200  23.300 10.500  24.000 10.500  24.000 
      12.500  23.300 12.500  23.300 20.600  23.500 20.600  23.500 25.200  
      22.100 25.200  22.100 20.600  22.300 20.600  22.300 12.500  22.000 
      12.500  22.000 11.500  17.300 11.500  17.300 20.600  17.500 20.600  
      17.500 25.200  16.100 25.200  16.100 20.600  16.300 20.600  16.300 
      11.500  11.300 11.500  11.300 20.600  11.500 20.600  11.500 25.200  
      10.100 25.200  10.100 20.600  10.300 20.600  10.300 11.500  5.300 11.500 
       5.300 20.600  5.500 20.600  5.500 25.200  4.100 25.200  ;
    LAYER ML2 ;
      POLYGON 22.000 12.500  22.000 10.500  24.000 10.500  24.000 12.500  
      22.000 12.500  ;
      POLYGON 1.000 14.500  1.000 16.500  3.000 16.500  3.000 14.500  1.000 
      14.500  ;
    LAYER POL ;
      POLYGON 1.000 16.500  1.000 14.500  2.800 14.500  2.800 1.700  3.800 
      1.700  3.800 14.500  5.800 14.500  5.800 1.700  6.800 1.700  6.800 
      14.500  8.800 14.500  8.800 1.700  9.800 1.700  9.800 14.500  11.800 
      14.500  11.800 1.700  12.800 1.700  12.800 14.500  14.800 14.500  14.800 
      1.700  15.800 1.700  15.800 14.500  17.800 14.500  17.800 1.700  18.800 
      1.700  18.800 14.500  20.800 14.500  20.800 1.700  21.800 1.700  21.800 
      14.500  23.800 14.500  23.800 1.700  24.800 1.700  24.800 26.500  23.800 
      26.500  23.800 16.500  21.800 16.500  21.800 26.500  20.800 26.500  
      20.800 16.500  18.800 16.500  18.800 26.500  17.800 26.500  17.800 
      16.500  15.800 16.500  15.800 26.500  14.800 26.500  14.800 16.500  
      12.800 16.500  12.800 26.500  11.800 26.500  11.800 16.500  9.800 16.500 
       9.800 26.500  8.800 26.500  8.800 16.500  6.800 16.500  6.800 26.500  
      5.800 26.500  5.800 16.500  3.800 16.500  3.800 26.500  2.800 26.500  
      2.800 16.500  1.000 16.500  ;
    LAYER VIA1 ;
      POLYGON 22.500 11.000  22.500 12.000  23.500 12.000  23.500 11.000  
      22.500 11.000  ;
      POLYGON 1.500 15.000  1.500 16.000  2.500 16.000  2.500 15.000  1.500 
      15.000  ;
  END
END inv8LEF


END LIBRARY
