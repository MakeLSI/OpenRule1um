VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO nr31
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 12.500 BY 30.000 ;
  SYMMETRY X Y ;
  SITE unit ;
 
  PIN A
    USE SIGNAL ;
    PORT
      LAYER ML1 ;
        POLYGON 1.000 14.500  1.000 16.500  3.000 16.500  3.000 14.500  1.000 
        14.500  ;
    END
    PORT
      LAYER ML2 ;
        POLYGON 1.000 14.500  1.000 16.500  3.000 16.500  3.000 14.500  1.000 
        14.500  ;
    END
  END A
  PIN B
    USE SIGNAL ;
    PORT
      LAYER ML2 ;
        POLYGON 4.000 11.500  4.000 13.500  6.000 13.500  6.000 11.500  4.000 
        11.500  ;
    END
    PORT
      LAYER ML1 ;
        POLYGON 4.000 11.500  4.000 13.500  6.000 13.500  6.000 11.500  4.000 
        11.500  ;
    END
  END B
  PIN C
    USE SIGNAL ;
    PORT
      LAYER ML1 ;
        POLYGON 7.000 12.000  7.000 14.000  9.000 14.000  9.000 12.000  7.000 
        12.000  ;
    END
    PORT
      LAYER ML2 ;
        POLYGON 7.000 12.000  7.000 14.000  9.000 14.000  9.000 12.000  7.000 
        12.000  ;
    END
  END C
  PIN VDD
    USE POWER ;
    PORT
      LAYER ML1 ;
        RECT -0.500 28.500  13.000 30.500  ;
    END
  END VDD
  PIN VSS
    USE GROUND ;
    PORT
      LAYER ML1 ;
        RECT -0.500 -0.500  13.000 1.500  ;
    END
  END VSS

  PIN YB
    USE SIGNAL ;
    PORT
      LAYER ML1 ;
        RECT 10.000 7.800  12.000 9.800  ;
    END
    PORT
      LAYER ML2 ;
        RECT 10.000 7.800  12.000 9.800  ;
    END
    PORT
      LAYER ML1 ;
        WIDTH 1.000  ;
        PATH 4.800 3.800 4.800 6.300 10.800 6.300  ;
    END
    PORT
      LAYER ML1 ;
        WIDTH 1.000  ;
        PATH 9.800 20.500 9.800 18.000 10.800 18.000 10.800 3.800  ;
    END
  END YB
  OBS

    LAYER ML1 ;
      WIDTH 1.000  ;
      PATH 1.800 1.000 1.800 3.800  ;

      WIDTH 1.400  ;
      PATH 2.800 21.300 2.800 28.500  ;


      WIDTH 1.000  ;
      PATH 7.800 1.000 7.800 3.800  ;
      WIDTH 1.000  ;
      PATH 4.800 3.800 4.800 6.300 10.800 6.300  ;

      WIDTH 1.400  ;
      PATH 9.800 21.300 9.800 24.500  ;
      WIDTH 1.000  ;
      PATH 9.800 20.500 9.800 18.000 10.800 18.000 10.800 3.800  ;

    VIA 1.800 3.800  dcont ;
    VIA 2.800 22.500  dcont ;
    VIA 2.800 20.500  dcont ;
    VIA 2.800 24.500  dcont ;
    VIA 4.800 3.800  dcont ;
    VIA 7.800 3.800  dcont ;
    VIA 10.800 3.800  dcont ;
    VIA 9.800 20.500  dcont ;
    VIA 9.800 22.500  dcont ;
    VIA 9.800 24.500  dcont ;
    VIA 5.000 12.500  pcont ;
    VIA 8.200 29.500  nsubcont ;
    VIA 8.000 13.000  pcont ;
    VIA 2.000 15.500  pcont ;
    VIA 6.500 0.500  psubcont ;
  END
END nr31

MACRO dcont
  CLASS CORE ;
  OBS
    LAYER ML1 ;
      RECT -1.000 -1.000  1.000 1.000  ;
  END
END dcont

MACRO pcont
  CLASS CORE ;
  OBS
    LAYER ML1 ;
      RECT -1.000 -1.000  1.000 1.000  ;
  END
END pcont

MACRO nsubcont
  CLASS CORE ;
  OBS
    LAYER ML1 ;
      RECT -1.000 -1.000  1.000 1.000  ;
  END
END nsubcont

MACRO psubcont
  CLASS CORE ;
  OBS
    LAYER ML1 ;
      RECT -1.000 -1.000  1.000 1.000  ;
  END
END psubcont


END LIBRARY
