*******************************************************************************
* CDL netlist
*
* Library : OpenRule1um_StdCell
* Top Cell Name: sff1m2_r
* View Name: extracted
* Netlist created: 07.4.2020 15:22:50
*******************************************************************************

*.SCALE METER
*.GLOBAL VDD VSS

*******************************************************************************
* Library Name: OpenRule1um_StdCell
* Cell Name:    sff1m2_r
* View Name:    extracted
*******************************************************************************

.SUBCKT sff1m2_r

MM194 n4 n6 n2 n2 pch w=6e-06 l=1e-06 as=1.2e-11 ps=1e-05 ad=1.2e-11 pd=1e-05 $X=5.58e-05 $Y=2.08e-05
MM169 n1 n5 n16 n1 nch w=2e-06 l=1e-06 as=1e-12 ps=4e-06 ad=2e-12 pd=6e-06 $X=2.88e-05 $Y=2.8e-06
MM165 n1 n10 n14 n1 nch w=2e-06 l=1e-06 as=2e-12 ps=4e-06 ad=4e-12 pd=6e-06 $X=1.88e-05 $Y=2.8e-06
MM162 n1 n13 n12 n1 nch w=2e-06 l=1e-06 as=4e-12 ps=6e-06 ad=4e-12 pd=6e-06 $X=2.8e-06 $Y=2.8e-06
MM173 n0 n7 n18 n1 nch w=2e-06 l=1e-06 as=1e-12 ps=4e-06 ad=2e-12 pd=6e-06 $X=4.23e-05 $Y=2.8e-06
MM189 n22 n7 n0 n2 pch w=6e-06 l=1e-06 as=6e-12 ps=1e-05 ad=3e-12 pd=8e-06 $X=3.68e-05 $Y=2.08e-05
MM193 n6 n3 n2 n2 pch w=6e-06 l=1e-06 as=6e-12 ps=1e-05 ad=6e-12 pd=1e-05 $X=4.78e-05 $Y=2.08e-05
MM184 n5 n7 n21 n2 pch w=6e-06 l=1e-06 as=3e-12 ps=8e-06 ad=6e-12 pd=1e-05 $X=2.38e-05 $Y=2.08e-05
MM176 n19 n3 n6 n1 nch w=2e-06 l=1e-06 as=2e-12 ps=6e-06 ad=1e-12 pd=4e-06 $X=4.93e-05 $Y=2.8e-06
MM177 n4 n6 n1 n1 nch w=2e-06 l=1e-06 as=4e-12 ps=6e-06 ad=4e-12 pd=6e-06 $X=5.58e-05 $Y=2.8e-06
MM172 n17 n9 n0 n1 nch w=2e-06 l=1e-06 as=2e-12 ps=6e-06 ad=1e-12 pd=4e-06 $X=3.93e-05 $Y=2.8e-06
MM195 n2 n4 n8 n2 pch w=6e-06 l=1e-06 as=6e-12 ps=1e-05 ad=6e-12 pd=1e-05 $X=5.88e-05 $Y=2.08e-05
MM175 n1 n0 n19 n1 nch w=2e-06 l=1e-06 as=1e-12 ps=4e-06 ad=2e-12 pd=6e-06 $X=4.73e-05 $Y=2.8e-06
MM180 n9 n12 n2 n2 pch w=6e-06 l=1e-06 as=1.2e-11 ps=1e-05 ad=1.2e-11 pd=1e-05 $X=9.3e-06 $Y=2.08e-05
MM179 n2 n13 n12 n2 pch w=6e-06 l=1e-06 as=1.2e-11 ps=1e-05 ad=1.2e-11 pd=1e-05 $X=2.8e-06 $Y=1.95e-05
MM181 n2 n9 n7 n2 pch w=6e-06 l=1e-06 as=6e-12 ps=1e-05 ad=6e-12 pd=1e-05 $X=1.23e-05 $Y=2.08e-05
MM178 n1 n4 n8 n1 nch w=2e-06 l=1e-06 as=2e-12 ps=6e-06 ad=2e-12 pd=6e-06 $X=5.88e-05 $Y=2.8e-06
MM167 n5 n9 n15 n1 nch w=2e-06 l=1e-06 as=1e-12 ps=4e-06 ad=2e-12 pd=6e-06 $X=2.38e-05 $Y=2.8e-06
MM192 n2 n0 n6 n2 pch w=6e-06 l=1e-06 as=6e-12 ps=1e-05 ad=6e-12 pd=1e-05 $X=4.48e-05 $Y=2.08e-05
MM191 n23 n6 n2 n2 pch w=6e-06 l=1e-06 as=6e-12 ps=1e-05 ad=3e-12 pd=8e-06 $X=4.18e-05 $Y=2.08e-05
MM174 n18 n6 n1 n1 nch w=2e-06 l=1e-06 as=2e-12 ps=6e-06 ad=1e-12 pd=4e-06 $X=4.43e-05 $Y=2.8e-06
MM171 n1 n11 n17 n1 nch w=2e-06 l=1e-06 as=2e-12 ps=4e-06 ad=4e-12 pd=6e-06 $X=3.73e-05 $Y=2.8e-06
MM187 n11 n3 n2 n2 pch w=6e-06 l=1e-06 as=6e-12 ps=1e-05 ad=6e-12 pd=1e-05 $X=3.18e-05 $Y=2.08e-05
MM163 n9 n12 n1 n1 nch w=2e-06 l=1e-06 as=4e-12 ps=6e-06 ad=4e-12 pd=6e-06 $X=9.3e-06 $Y=2.8e-06
MM186 n2 n5 n11 n2 pch w=6e-06 l=1e-06 as=6e-12 ps=1e-05 ad=6e-12 pd=1e-05 $X=2.88e-05 $Y=2.08e-05
MM190 n0 n9 n23 n2 pch w=6e-06 l=1e-06 as=3e-12 ps=8e-06 ad=6e-12 pd=1e-05 $X=3.98e-05 $Y=2.08e-05
MM185 n21 n11 n2 n2 pch w=6e-06 l=1e-06 as=6e-12 ps=1e-05 ad=3e-12 pd=8e-06 $X=2.58e-05 $Y=2.08e-05
MM188 n2 n11 n22 n2 pch w=6e-06 l=1e-06 as=3e-12 ps=8e-06 ad=6e-12 pd=1e-05 $X=3.48e-05 $Y=2.08e-05
MM168 n15 n11 n1 n1 nch w=2e-06 l=1e-06 as=2e-12 ps=6e-06 ad=1e-12 pd=4e-06 $X=2.58e-05 $Y=2.8e-06
MM182 n2 n10 n20 n2 pch w=6e-06 l=1e-06 as=6e-12 ps=8e-06 ad=1.2e-11 pd=1e-05 $X=1.88e-05 $Y=2.08e-05
MM170 n16 n3 n11 n1 nch w=2e-06 l=1e-06 as=2e-12 ps=6e-06 ad=1e-12 pd=4e-06 $X=3.08e-05 $Y=2.8e-06
MM164 n1 n9 n7 n1 nch w=2e-06 l=1e-06 as=2e-12 ps=6e-06 ad=2e-12 pd=6e-06 $X=1.23e-05 $Y=2.8e-06
MM183 n20 n9 n5 n2 pch w=6e-06 l=1e-06 as=6e-12 ps=1e-05 ad=3e-12 pd=8e-06 $X=2.08e-05 $Y=2.08e-05
MM166 n14 n7 n5 n1 nch w=2e-06 l=1e-06 as=2e-12 ps=6e-06 ad=1e-12 pd=4e-06 $X=2.08e-05 $Y=2.8e-06
.ENDS
