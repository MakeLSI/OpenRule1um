*******************************************************************************
* CDL netlist
*
* Library : OpenRule1um_StdCell
* Top Cell Name: sff1_r
* View Name: extracted
* Netlist created: 07.4.2020 15:15:01
*******************************************************************************

*.SCALE METER
*.GLOBAL VDD VSS

*******************************************************************************
* Library Name: OpenRule1um_StdCell
* Cell Name:    sff1_r
* View Name:    extracted
*******************************************************************************

.SUBCKT sff1_r

MM146 n9 n12 n2 n2 pch w=6e-06 l=1e-06 as=1.2e-11 ps=1e-05 ad=1.2e-11 pd=1e-05 $X=9.3e-06 $Y=2.08e-05
MM130 n1 n9 n8 n1 nch w=2e-06 l=1e-06 as=2e-12 ps=6e-06 ad=2e-12 pd=6e-06 $X=1.23e-05 $Y=2.8e-06
MM140 n18 n7 n1 n1 nch w=2e-06 l=1e-06 as=2e-12 ps=6e-06 ad=1e-12 pd=4e-06 $X=4.43e-05 $Y=2.8e-06
MM139 n0 n8 n18 n1 nch w=2e-06 l=1e-06 as=1e-12 ps=4e-06 ad=2e-12 pd=6e-06 $X=4.23e-05 $Y=2.8e-06
MM147 n2 n9 n8 n2 pch w=6e-06 l=1e-06 as=6e-12 ps=1e-05 ad=6e-12 pd=1e-05 $X=1.23e-05 $Y=2.08e-05
MM138 n17 n9 n0 n1 nch w=2e-06 l=1e-06 as=2e-12 ps=6e-06 ad=1e-12 pd=4e-06 $X=3.93e-05 $Y=2.8e-06
MM159 n7 n5 n2 n2 pch w=6e-06 l=1e-06 as=6e-12 ps=1e-05 ad=6e-12 pd=1e-05 $X=4.93e-05 $Y=2.08e-05
MM153 n3 n5 n2 n2 pch w=6e-06 l=1e-06 as=6e-12 ps=1e-05 ad=6e-12 pd=1e-05 $X=3.18e-05 $Y=2.08e-05
MM161 n2 n4 n11 n2 pch w=6e-06 l=1e-06 as=6e-12 ps=1e-05 ad=6e-12 pd=1e-05 $X=5.88e-05 $Y=2.08e-05
MM160 n4 n7 n2 n2 pch w=6e-06 l=1e-06 as=1.2e-11 ps=1e-05 ad=1.2e-11 pd=1e-05 $X=5.58e-05 $Y=2.08e-05
MM151 n21 n3 n2 n2 pch w=6e-06 l=1e-06 as=6e-12 ps=1e-05 ad=3e-12 pd=8e-06 $X=2.58e-05 $Y=2.08e-05
MM156 n0 n9 n23 n2 pch w=6e-06 l=1e-06 as=3e-12 ps=8e-06 ad=6e-12 pd=1e-05 $X=4.13e-05 $Y=2.08e-05
MM144 n1 n4 n11 n1 nch w=2e-06 l=1e-06 as=2e-12 ps=6e-06 ad=2e-12 pd=6e-06 $X=5.88e-05 $Y=2.8e-06
MM148 n2 n10 n20 n2 pch w=6e-06 l=1e-06 as=6e-12 ps=8e-06 ad=1.2e-11 pd=1e-05 $X=1.88e-05 $Y=2.08e-05
MM143 n4 n7 n1 n1 nch w=2e-06 l=1e-06 as=4e-12 ps=6e-06 ad=4e-12 pd=6e-06 $X=5.58e-05 $Y=2.8e-06
MM134 n15 n3 n1 n1 nch w=2e-06 l=1e-06 as=2e-12 ps=6e-06 ad=1e-12 pd=4e-06 $X=2.58e-05 $Y=2.8e-06
MM142 n19 n5 n7 n1 nch w=2e-06 l=1e-06 as=2e-12 ps=6e-06 ad=1e-12 pd=4e-06 $X=4.93e-05 $Y=2.8e-06
MM132 n14 n8 n6 n1 nch w=2e-06 l=1e-06 as=2e-12 ps=6e-06 ad=1e-12 pd=4e-06 $X=2.08e-05 $Y=2.8e-06
MM145 n2 n13 n12 n2 pch w=6e-06 l=1e-06 as=1.2e-11 ps=1e-05 ad=1.2e-11 pd=1e-05 $X=2.8e-06 $Y=1.95e-05
MM129 n9 n12 n1 n1 nch w=2e-06 l=1e-06 as=4e-12 ps=6e-06 ad=4e-12 pd=6e-06 $X=9.3e-06 $Y=2.8e-06
MM158 n2 n0 n7 n2 pch w=6e-06 l=1e-06 as=6e-12 ps=1e-05 ad=6e-12 pd=1e-05 $X=4.63e-05 $Y=2.08e-05
MM157 n23 n7 n2 n2 pch w=6e-06 l=1e-06 as=6e-12 ps=1e-05 ad=3e-12 pd=8e-06 $X=4.33e-05 $Y=2.08e-05
MM131 n1 n10 n14 n1 nch w=2e-06 l=1e-06 as=2e-12 ps=4e-06 ad=4e-12 pd=6e-06 $X=1.88e-05 $Y=2.8e-06
MM128 n1 n13 n12 n1 nch w=2e-06 l=1e-06 as=4e-12 ps=6e-06 ad=4e-12 pd=6e-06 $X=2.8e-06 $Y=2.8e-06
MM155 n22 n8 n0 n2 pch w=6e-06 l=1e-06 as=6e-12 ps=1e-05 ad=7.5e-12 pd=1.1e-05 $X=3.83e-05 $Y=2.08e-05
MM150 n6 n8 n21 n2 pch w=6e-06 l=1e-06 as=3e-12 ps=8e-06 ad=6e-12 pd=1e-05 $X=2.38e-05 $Y=2.08e-05
MM141 n1 n0 n19 n1 nch w=2e-06 l=1e-06 as=1e-12 ps=4e-06 ad=2e-12 pd=6e-06 $X=4.73e-05 $Y=2.8e-06
MM135 n1 n6 n16 n1 nch w=2e-06 l=1e-06 as=1e-12 ps=4e-06 ad=2e-12 pd=6e-06 $X=2.88e-05 $Y=2.8e-06
MM137 n1 n3 n17 n1 nch w=2e-06 l=1e-06 as=2e-12 ps=4e-06 ad=4e-12 pd=6e-06 $X=3.73e-05 $Y=2.8e-06
MM154 n2 n3 n22 n2 pch w=6e-06 l=1e-06 as=7.5e-12 ps=1.1e-05 ad=6e-12 pd=1e-05 $X=3.48e-05 $Y=2.08e-05
MM149 n20 n9 n6 n2 pch w=6e-06 l=1e-06 as=6e-12 ps=1e-05 ad=3e-12 pd=8e-06 $X=2.08e-05 $Y=2.08e-05
MM133 n6 n9 n15 n1 nch w=2e-06 l=1e-06 as=1e-12 ps=4e-06 ad=2e-12 pd=6e-06 $X=2.38e-05 $Y=2.8e-06
MM136 n16 n5 n3 n1 nch w=2e-06 l=1e-06 as=2e-12 ps=6e-06 ad=1e-12 pd=4e-06 $X=3.08e-05 $Y=2.8e-06
MM152 n2 n6 n3 n2 pch w=6e-06 l=1e-06 as=6e-12 ps=1e-05 ad=6e-12 pd=1e-05 $X=2.88e-05 $Y=2.08e-05
.ENDS
