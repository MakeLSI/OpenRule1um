VERSION 5.3 ;

NAMESCASESENSITIVE ON ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS











MACRO nr21LEF
  CLASS BLOCK ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER POL ;
        POLYGON 1.000 16.500  1.000 14.500  2.000 14.500  2.000 9.500  2.800 
        9.500  2.800 1.700  3.800 1.700  3.800 10.500  3.000 10.500  3.000 
        17.100  4.300 17.100  4.300 26.500  3.300 26.500  3.300 18.100  2.000 
        18.100  2.000 16.500  1.000 16.500  ;
    END
    PORT
      LAYER ML1 ;
        POLYGON 1.000 14.500  1.000 16.500  3.000 16.500  3.000 14.500  1.000 
        14.500  ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER POL ;
        POLYGON 4.000 13.500  4.000 11.500  5.000 11.500  5.000 9.500  5.800 
        9.500  5.800 1.700  6.800 1.700  6.800 10.500  6.000 10.500  6.000 
        15.000  6.300 15.000  6.300 26.500  5.300 26.500  5.300 16.000  5.000 
        16.000  5.000 13.500  4.000 13.500  ;
    END
    PORT
      LAYER ML1 ;
        POLYGON 4.000 11.500  4.000 13.500  6.000 13.500  6.000 11.500  4.000 
        11.500  ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    PORT
      LAYER ML1 ;
        POLYGON -0.500 30.500  -0.500 28.500  1.600 28.500  1.600 20.600  
        3.000 20.600  3.000 28.500  10.000 28.500  10.000 30.500  -0.500 
        30.500  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    PORT
      LAYER ML1 ;
        POLYGON -0.500 1.500  -0.500 -0.500  10.000 -0.500  10.000 1.500  
        8.300 1.500  8.300 4.200  7.300 4.200  7.300 1.500  2.300 1.500  2.300 
        4.200  1.300 4.200  1.300 1.500  -0.500 1.500  ;
    END
  END VSS
  PIN YB
    DIRECTION OUTPUT ;
    PORT
      LAYER ML1 ;
        POLYGON 4.300 6.700  4.300 3.200  5.300 3.200  5.300 5.700  8.300 
        5.700  8.300 8.500  9.000 8.500  9.000 10.500  8.300 10.500  8.300 
        16.000  7.800 16.000  7.800 20.600  8.000 20.600  8.000 25.200  6.600 
        25.200  6.600 20.600  6.800 20.600  6.800 15.000  7.300 15.000  7.300 
        10.500  7.000 10.500  7.000 8.500  7.300 8.500  7.300 6.700  4.300 
        6.700  ;
    END
  END YB
  OBS
    LAYER CNT ;
      POLYGON 1.800 20.000  1.800 21.000  2.800 21.000  2.800 20.000  1.800 
      20.000  ;
      POLYGON 1.800 24.000  1.800 25.000  2.800 25.000  2.800 24.000  1.800 
      24.000  ;
      POLYGON 4.300 3.200  4.300 4.200  5.300 4.200  5.300 3.200  4.300 3.200  ;
      
      POLYGON 7.300 3.200  7.300 4.200  8.300 4.200  8.300 3.200  7.300 3.200  ;
      
      POLYGON 6.800 20.000  6.800 21.000  7.800 21.000  7.800 20.000  6.800 
      20.000  ;
      POLYGON 6.800 22.000  6.800 23.000  7.800 23.000  7.800 22.000  6.800 
      22.000  ;
      POLYGON 6.800 24.000  6.800 25.000  7.800 25.000  7.800 24.000  6.800 
      24.000  ;
      POLYGON 4.500 12.000  4.500 13.000  5.500 13.000  5.500 12.000  4.500 
      12.000  ;
      POLYGON 5.000 29.000  5.000 30.000  6.000 30.000  6.000 29.000  5.000 
      29.000  ;
      POLYGON 1.500 15.000  1.500 16.000  2.500 16.000  2.500 15.000  1.500 
      15.000  ;
      POLYGON 4.500 0.000  4.500 1.000  5.500 1.000  5.500 0.000  4.500 0.000  ;
      
      POLYGON 1.800 22.000  1.800 23.000  2.800 23.000  2.800 22.000  1.800 
      22.000  ;
      POLYGON 1.300 3.200  1.300 4.200  2.300 4.200  2.300 3.200  1.300 3.200  ;
      
    LAYER FRAME ;
      POLYGON 0.000 0.000  9.500 0.000  9.500 30.000  0.000 30.000  0.000 
      0.000  ;
      RECT -0.500 -0.500  10.000 1.500  ;
      RECT -0.500 28.500  10.000 30.500  ;
    LAYER ML1 ;
      POLYGON 4.000 11.500  4.000 13.500  6.000 13.500  6.000 11.500  4.000 
      11.500  ;
      RECT 4.000 -0.500  6.000 1.500  ;
      POLYGON 1.000 14.500  1.000 16.500  3.000 16.500  3.000 14.500  1.000 
      14.500  ;
      RECT 1.000 14.500  3.000 16.500  ;
      RECT 4.500 28.500  6.500 30.500  ;
      RECT 4.000 11.500  6.000 13.500  ;
      RECT 6.300 23.500  8.300 25.500  ;
      RECT 6.300 21.500  8.300 23.500  ;
      RECT 6.300 19.500  8.300 21.500  ;
      RECT 6.800 2.700  8.800 4.700  ;
      RECT 3.800 2.700  5.800 4.700  ;
      RECT 1.300 23.500  3.300 25.500  ;
      RECT 1.300 19.500  3.300 21.500  ;
      RECT 1.300 21.500  3.300 23.500  ;
      RECT 0.800 2.700  2.800 4.700  ;
      POLYGON -0.500 30.500  -0.500 28.500  1.600 28.500  1.600 20.600  3.000 
      20.600  3.000 28.500  10.000 28.500  10.000 30.500  -0.500 30.500  ;
      POLYGON -0.500 1.500  -0.500 -0.500  10.000 -0.500  10.000 1.500  8.300 
      1.500  8.300 4.200  7.300 4.200  7.300 1.500  2.300 1.500  2.300 4.200  
      1.300 4.200  1.300 1.500  -0.500 1.500  ;
      POLYGON 4.300 6.700  4.300 3.200  5.300 3.200  5.300 5.700  8.300 5.700  
      8.300 8.500  9.000 8.500  9.000 10.500  8.300 10.500  8.300 16.000  
      7.800 16.000  7.800 20.600  8.000 20.600  8.000 25.200  6.600 25.200  
      6.600 20.600  6.800 20.600  6.800 15.000  7.300 15.000  7.300 10.500  
      7.000 10.500  7.000 8.500  7.300 8.500  7.300 6.700  4.300 6.700  ;
    LAYER ML2 ;
      POLYGON 4.000 11.500  4.000 13.500  6.000 13.500  6.000 11.500  4.000 
      11.500  ;
      POLYGON 7.000 8.500  7.000 10.500  9.000 10.500  9.000 8.500  7.000 
      8.500  ;
      POLYGON 1.000 14.500  1.000 16.500  3.000 16.500  3.000 14.500  1.000 
      14.500  ;
    LAYER POL ;
      POLYGON 4.000 13.500  4.000 11.500  5.000 11.500  5.000 9.500  5.800 
      9.500  5.800 1.700  6.800 1.700  6.800 10.500  6.000 10.500  6.000 
      15.000  6.300 15.000  6.300 26.500  5.300 26.500  5.300 16.000  5.000 
      16.000  5.000 13.500  4.000 13.500  ;
      POLYGON 1.000 16.500  1.000 14.500  2.000 14.500  2.000 9.500  2.800 
      9.500  2.800 1.700  3.800 1.700  3.800 10.500  3.000 10.500  3.000 
      17.100  4.300 17.100  4.300 26.500  3.300 26.500  3.300 18.100  2.000 
      18.100  2.000 16.500  1.000 16.500  ;
    LAYER VIA1 ;
      POLYGON 4.500 12.000  4.500 13.000  5.500 13.000  5.500 12.000  4.500 
      12.000  ;
      POLYGON 7.500 9.000  7.500 10.000  8.500 10.000  8.500 9.000  7.500 
      9.000  ;
      POLYGON 1.500 15.000  1.500 16.000  2.500 16.000  2.500 15.000  1.500 
      15.000  ;
  END
END nr21LEF


END LIBRARY
