VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO na41
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 15.500 BY 30.000 ;
  SYMMETRY X Y ;
  SITE unit ;
 
  PIN A
    USE SIGNAL ;
    PORT
      LAYER ML2 ;
        POLYGON 1.000 15.500  1.000 17.500  3.000 17.500  3.000 15.500  1.000 
        15.500  ;
    END
    PORT
      LAYER ML1 ;
        POLYGON 1.000 15.500  1.000 17.500  3.000 17.500  3.000 15.500  1.000 
        15.500  ;
    END
  END A
  PIN B
    USE SIGNAL ;
    PORT
      LAYER ML2 ;
        POLYGON 4.000 12.500  4.000 14.500  6.000 14.500  6.000 12.500  4.000 
        12.500  ;
    END
    PORT
      LAYER ML1 ;
        POLYGON 4.000 12.500  4.000 14.500  6.000 14.500  6.000 12.500  4.000 
        12.500  ;
    END
  END B
  PIN C
    USE SIGNAL ;
    PORT
      LAYER ML2 ;
        POLYGON 7.000 9.500  7.000 11.500  9.000 11.500  9.000 9.500  7.000 
        9.500  ;
    END
    PORT
      LAYER ML1 ;
        POLYGON 7.000 9.500  7.000 11.500  9.000 11.500  9.000 9.500  7.000 
        9.500  ;
    END
  END C
  PIN D
    USE SIGNAL ;
    PORT
      LAYER ML2 ;
        POLYGON 10.000 6.500  10.000 8.500  12.000 8.500  12.000 6.500  10.000 
        6.500  ;
    END
    PORT
      LAYER ML1 ;
        POLYGON 10.000 6.500  10.000 8.500  12.000 8.500  12.000 6.500  10.000 
        6.500  ;
    END
  END D
  PIN VDD
    USE POWER ;
    PORT
      LAYER ML1 ;
        RECT -0.500 28.500  16.000 30.500  ;
    END
  END VDD
  PIN VSS
    USE GROUND ;
    PORT
      LAYER ML1 ;
        RECT -0.500 -0.500  16.000 1.500  ;
    END
  END VSS
  PIN YB
    USE SIGNAL ;
    PORT
      LAYER ML1 ;
        POLYGON 13.000 9.500  13.000 11.500  15.000 11.500  15.000 9.500  
        13.000 9.500  ;
    END
    PORT
      LAYER ML2 ;
        POLYGON 13.000 9.500  13.000 11.500  15.000 11.500  15.000 9.500  
        13.000 9.500  ;
    END
    PORT
      LAYER ML1 ;
        WIDTH 1.000  ;
        PATH 10.800 20.500 10.800 18.000  ;
    END
    PORT
      LAYER ML1 ;
        WIDTH 1.000  ;
        PATH 4.800 20.500 4.800 18.000 13.800 18.000 13.800 3.800 10.800 3.800 
         ;
    END
  END YB
  OBS

    LAYER ML1 ;
      WIDTH 1.400  ;
      PATH 1.800 21.300 1.800 28.500  ;
      WIDTH 1.000  ;
      PATH 1.800 1.000 1.800 3.800  ;
      WIDTH 1.400  ;
      PATH 4.800 21.300 4.800 24.500  ;

      WIDTH 1.400  ;
      PATH 7.800 21.300 7.800 28.500  ;
      WIDTH 1.000  ;
      PATH 4.800 20.500 4.800 18.000 13.800 18.000 13.800 3.800 10.800 3.800 
       ;
      WIDTH 1.000  ;
      PATH 10.800 20.500 10.800 18.000  ;
      WIDTH 1.400  ;
      PATH 10.800 21.300 10.800 24.500  ;
      WIDTH 1.400  ;
      PATH 13.800 21.300 13.800 28.500  ;
      WIDTH 1.400  ;
      PATH 13.800 21.300 13.800 24.500  ;

    VIA 1.800 22.500  dcont ;
    VIA 1.800 20.500  dcont ;
    VIA 1.800 3.800  dcont ;
    VIA 1.800 24.500  dcont ;
    VIA 4.800 22.500  dcont ;
    VIA 4.800 20.500  dcont ;
    VIA 4.800 24.500  dcont ;
    VIA 7.800 24.500  dcont ;
    VIA 7.800 22.500  dcont ;
    VIA 7.800 20.500  dcont ;
    VIA 10.800 3.800  dcont ;
    VIA 10.800 20.500  dcont ;
    VIA 10.800 22.500  dcont ;
    VIA 10.800 24.500  dcont ;
    VIA 13.800 24.500  dcont ;
    VIA 13.800 22.500  dcont ;
    VIA 13.800 20.500  dcont ;
    VIA 11.000 7.500  pcont ;
    VIA 8.000 10.500  pcont ;
    VIA 5.500 29.500  nsubcont ;
    VIA 5.000 13.500  pcont ;
    VIA 2.000 16.500  pcont ;
    VIA 5.000 0.500  psubcont ;
  END
END na41

MACRO dcont
  CLASS CORE ;
  OBS
    LAYER ML1 ;
      RECT -1.000 -1.000  1.000 1.000  ;
  END
END dcont

MACRO pcont
  CLASS CORE ;
  OBS
    LAYER ML1 ;
      RECT -1.000 -1.000  1.000 1.000  ;
  END
END pcont

MACRO nsubcont
  CLASS CORE ;
  OBS
    LAYER ML1 ;
      RECT -1.000 -1.000  1.000 1.000  ;
  END
END nsubcont

MACRO psubcont
  CLASS CORE ;
  OBS
    LAYER ML1 ;
      RECT -1.000 -1.000  1.000 1.000  ;
  END
END psubcont


END LIBRARY
